module ShiftRegister2034(
    input data_in,
    output [2033:0] data_out,
    input clock,
    input enable,
    input nreset
);
    reg [2033:0] r_data;
    always @(posedge clock) begin
        if (!nreset) begin
            r_data <= 0;
        end else begin
            if (enable) begin
                
                r_data[0] <= data_in;
                
                r_data[1] <= r_data[0];
                
                r_data[2] <= r_data[1];
                
                r_data[3] <= r_data[2];
                
                r_data[4] <= r_data[3];
                
                r_data[5] <= r_data[4];
                
                r_data[6] <= r_data[5];
                
                r_data[7] <= r_data[6];
                
                r_data[8] <= r_data[7];
                
                r_data[9] <= r_data[8];
                
                r_data[10] <= r_data[9];
                
                r_data[11] <= r_data[10];
                
                r_data[12] <= r_data[11];
                
                r_data[13] <= r_data[12];
                
                r_data[14] <= r_data[13];
                
                r_data[15] <= r_data[14];
                
                r_data[16] <= r_data[15];
                
                r_data[17] <= r_data[16];
                
                r_data[18] <= r_data[17];
                
                r_data[19] <= r_data[18];
                
                r_data[20] <= r_data[19];
                
                r_data[21] <= r_data[20];
                
                r_data[22] <= r_data[21];
                
                r_data[23] <= r_data[22];
                
                r_data[24] <= r_data[23];
                
                r_data[25] <= r_data[24];
                
                r_data[26] <= r_data[25];
                
                r_data[27] <= r_data[26];
                
                r_data[28] <= r_data[27];
                
                r_data[29] <= r_data[28];
                
                r_data[30] <= r_data[29];
                
                r_data[31] <= r_data[30];
                
                r_data[32] <= r_data[31];
                
                r_data[33] <= r_data[32];
                
                r_data[34] <= r_data[33];
                
                r_data[35] <= r_data[34];
                
                r_data[36] <= r_data[35];
                
                r_data[37] <= r_data[36];
                
                r_data[38] <= r_data[37];
                
                r_data[39] <= r_data[38];
                
                r_data[40] <= r_data[39];
                
                r_data[41] <= r_data[40];
                
                r_data[42] <= r_data[41];
                
                r_data[43] <= r_data[42];
                
                r_data[44] <= r_data[43];
                
                r_data[45] <= r_data[44];
                
                r_data[46] <= r_data[45];
                
                r_data[47] <= r_data[46];
                
                r_data[48] <= r_data[47];
                
                r_data[49] <= r_data[48];
                
                r_data[50] <= r_data[49];
                
                r_data[51] <= r_data[50];
                
                r_data[52] <= r_data[51];
                
                r_data[53] <= r_data[52];
                
                r_data[54] <= r_data[53];
                
                r_data[55] <= r_data[54];
                
                r_data[56] <= r_data[55];
                
                r_data[57] <= r_data[56];
                
                r_data[58] <= r_data[57];
                
                r_data[59] <= r_data[58];
                
                r_data[60] <= r_data[59];
                
                r_data[61] <= r_data[60];
                
                r_data[62] <= r_data[61];
                
                r_data[63] <= r_data[62];
                
                r_data[64] <= r_data[63];
                
                r_data[65] <= r_data[64];
                
                r_data[66] <= r_data[65];
                
                r_data[67] <= r_data[66];
                
                r_data[68] <= r_data[67];
                
                r_data[69] <= r_data[68];
                
                r_data[70] <= r_data[69];
                
                r_data[71] <= r_data[70];
                
                r_data[72] <= r_data[71];
                
                r_data[73] <= r_data[72];
                
                r_data[74] <= r_data[73];
                
                r_data[75] <= r_data[74];
                
                r_data[76] <= r_data[75];
                
                r_data[77] <= r_data[76];
                
                r_data[78] <= r_data[77];
                
                r_data[79] <= r_data[78];
                
                r_data[80] <= r_data[79];
                
                r_data[81] <= r_data[80];
                
                r_data[82] <= r_data[81];
                
                r_data[83] <= r_data[82];
                
                r_data[84] <= r_data[83];
                
                r_data[85] <= r_data[84];
                
                r_data[86] <= r_data[85];
                
                r_data[87] <= r_data[86];
                
                r_data[88] <= r_data[87];
                
                r_data[89] <= r_data[88];
                
                r_data[90] <= r_data[89];
                
                r_data[91] <= r_data[90];
                
                r_data[92] <= r_data[91];
                
                r_data[93] <= r_data[92];
                
                r_data[94] <= r_data[93];
                
                r_data[95] <= r_data[94];
                
                r_data[96] <= r_data[95];
                
                r_data[97] <= r_data[96];
                
                r_data[98] <= r_data[97];
                
                r_data[99] <= r_data[98];
                
                r_data[100] <= r_data[99];
                
                r_data[101] <= r_data[100];
                
                r_data[102] <= r_data[101];
                
                r_data[103] <= r_data[102];
                
                r_data[104] <= r_data[103];
                
                r_data[105] <= r_data[104];
                
                r_data[106] <= r_data[105];
                
                r_data[107] <= r_data[106];
                
                r_data[108] <= r_data[107];
                
                r_data[109] <= r_data[108];
                
                r_data[110] <= r_data[109];
                
                r_data[111] <= r_data[110];
                
                r_data[112] <= r_data[111];
                
                r_data[113] <= r_data[112];
                
                r_data[114] <= r_data[113];
                
                r_data[115] <= r_data[114];
                
                r_data[116] <= r_data[115];
                
                r_data[117] <= r_data[116];
                
                r_data[118] <= r_data[117];
                
                r_data[119] <= r_data[118];
                
                r_data[120] <= r_data[119];
                
                r_data[121] <= r_data[120];
                
                r_data[122] <= r_data[121];
                
                r_data[123] <= r_data[122];
                
                r_data[124] <= r_data[123];
                
                r_data[125] <= r_data[124];
                
                r_data[126] <= r_data[125];
                
                r_data[127] <= r_data[126];
                
                r_data[128] <= r_data[127];
                
                r_data[129] <= r_data[128];
                
                r_data[130] <= r_data[129];
                
                r_data[131] <= r_data[130];
                
                r_data[132] <= r_data[131];
                
                r_data[133] <= r_data[132];
                
                r_data[134] <= r_data[133];
                
                r_data[135] <= r_data[134];
                
                r_data[136] <= r_data[135];
                
                r_data[137] <= r_data[136];
                
                r_data[138] <= r_data[137];
                
                r_data[139] <= r_data[138];
                
                r_data[140] <= r_data[139];
                
                r_data[141] <= r_data[140];
                
                r_data[142] <= r_data[141];
                
                r_data[143] <= r_data[142];
                
                r_data[144] <= r_data[143];
                
                r_data[145] <= r_data[144];
                
                r_data[146] <= r_data[145];
                
                r_data[147] <= r_data[146];
                
                r_data[148] <= r_data[147];
                
                r_data[149] <= r_data[148];
                
                r_data[150] <= r_data[149];
                
                r_data[151] <= r_data[150];
                
                r_data[152] <= r_data[151];
                
                r_data[153] <= r_data[152];
                
                r_data[154] <= r_data[153];
                
                r_data[155] <= r_data[154];
                
                r_data[156] <= r_data[155];
                
                r_data[157] <= r_data[156];
                
                r_data[158] <= r_data[157];
                
                r_data[159] <= r_data[158];
                
                r_data[160] <= r_data[159];
                
                r_data[161] <= r_data[160];
                
                r_data[162] <= r_data[161];
                
                r_data[163] <= r_data[162];
                
                r_data[164] <= r_data[163];
                
                r_data[165] <= r_data[164];
                
                r_data[166] <= r_data[165];
                
                r_data[167] <= r_data[166];
                
                r_data[168] <= r_data[167];
                
                r_data[169] <= r_data[168];
                
                r_data[170] <= r_data[169];
                
                r_data[171] <= r_data[170];
                
                r_data[172] <= r_data[171];
                
                r_data[173] <= r_data[172];
                
                r_data[174] <= r_data[173];
                
                r_data[175] <= r_data[174];
                
                r_data[176] <= r_data[175];
                
                r_data[177] <= r_data[176];
                
                r_data[178] <= r_data[177];
                
                r_data[179] <= r_data[178];
                
                r_data[180] <= r_data[179];
                
                r_data[181] <= r_data[180];
                
                r_data[182] <= r_data[181];
                
                r_data[183] <= r_data[182];
                
                r_data[184] <= r_data[183];
                
                r_data[185] <= r_data[184];
                
                r_data[186] <= r_data[185];
                
                r_data[187] <= r_data[186];
                
                r_data[188] <= r_data[187];
                
                r_data[189] <= r_data[188];
                
                r_data[190] <= r_data[189];
                
                r_data[191] <= r_data[190];
                
                r_data[192] <= r_data[191];
                
                r_data[193] <= r_data[192];
                
                r_data[194] <= r_data[193];
                
                r_data[195] <= r_data[194];
                
                r_data[196] <= r_data[195];
                
                r_data[197] <= r_data[196];
                
                r_data[198] <= r_data[197];
                
                r_data[199] <= r_data[198];
                
                r_data[200] <= r_data[199];
                
                r_data[201] <= r_data[200];
                
                r_data[202] <= r_data[201];
                
                r_data[203] <= r_data[202];
                
                r_data[204] <= r_data[203];
                
                r_data[205] <= r_data[204];
                
                r_data[206] <= r_data[205];
                
                r_data[207] <= r_data[206];
                
                r_data[208] <= r_data[207];
                
                r_data[209] <= r_data[208];
                
                r_data[210] <= r_data[209];
                
                r_data[211] <= r_data[210];
                
                r_data[212] <= r_data[211];
                
                r_data[213] <= r_data[212];
                
                r_data[214] <= r_data[213];
                
                r_data[215] <= r_data[214];
                
                r_data[216] <= r_data[215];
                
                r_data[217] <= r_data[216];
                
                r_data[218] <= r_data[217];
                
                r_data[219] <= r_data[218];
                
                r_data[220] <= r_data[219];
                
                r_data[221] <= r_data[220];
                
                r_data[222] <= r_data[221];
                
                r_data[223] <= r_data[222];
                
                r_data[224] <= r_data[223];
                
                r_data[225] <= r_data[224];
                
                r_data[226] <= r_data[225];
                
                r_data[227] <= r_data[226];
                
                r_data[228] <= r_data[227];
                
                r_data[229] <= r_data[228];
                
                r_data[230] <= r_data[229];
                
                r_data[231] <= r_data[230];
                
                r_data[232] <= r_data[231];
                
                r_data[233] <= r_data[232];
                
                r_data[234] <= r_data[233];
                
                r_data[235] <= r_data[234];
                
                r_data[236] <= r_data[235];
                
                r_data[237] <= r_data[236];
                
                r_data[238] <= r_data[237];
                
                r_data[239] <= r_data[238];
                
                r_data[240] <= r_data[239];
                
                r_data[241] <= r_data[240];
                
                r_data[242] <= r_data[241];
                
                r_data[243] <= r_data[242];
                
                r_data[244] <= r_data[243];
                
                r_data[245] <= r_data[244];
                
                r_data[246] <= r_data[245];
                
                r_data[247] <= r_data[246];
                
                r_data[248] <= r_data[247];
                
                r_data[249] <= r_data[248];
                
                r_data[250] <= r_data[249];
                
                r_data[251] <= r_data[250];
                
                r_data[252] <= r_data[251];
                
                r_data[253] <= r_data[252];
                
                r_data[254] <= r_data[253];
                
                r_data[255] <= r_data[254];
                
                r_data[256] <= r_data[255];
                
                r_data[257] <= r_data[256];
                
                r_data[258] <= r_data[257];
                
                r_data[259] <= r_data[258];
                
                r_data[260] <= r_data[259];
                
                r_data[261] <= r_data[260];
                
                r_data[262] <= r_data[261];
                
                r_data[263] <= r_data[262];
                
                r_data[264] <= r_data[263];
                
                r_data[265] <= r_data[264];
                
                r_data[266] <= r_data[265];
                
                r_data[267] <= r_data[266];
                
                r_data[268] <= r_data[267];
                
                r_data[269] <= r_data[268];
                
                r_data[270] <= r_data[269];
                
                r_data[271] <= r_data[270];
                
                r_data[272] <= r_data[271];
                
                r_data[273] <= r_data[272];
                
                r_data[274] <= r_data[273];
                
                r_data[275] <= r_data[274];
                
                r_data[276] <= r_data[275];
                
                r_data[277] <= r_data[276];
                
                r_data[278] <= r_data[277];
                
                r_data[279] <= r_data[278];
                
                r_data[280] <= r_data[279];
                
                r_data[281] <= r_data[280];
                
                r_data[282] <= r_data[281];
                
                r_data[283] <= r_data[282];
                
                r_data[284] <= r_data[283];
                
                r_data[285] <= r_data[284];
                
                r_data[286] <= r_data[285];
                
                r_data[287] <= r_data[286];
                
                r_data[288] <= r_data[287];
                
                r_data[289] <= r_data[288];
                
                r_data[290] <= r_data[289];
                
                r_data[291] <= r_data[290];
                
                r_data[292] <= r_data[291];
                
                r_data[293] <= r_data[292];
                
                r_data[294] <= r_data[293];
                
                r_data[295] <= r_data[294];
                
                r_data[296] <= r_data[295];
                
                r_data[297] <= r_data[296];
                
                r_data[298] <= r_data[297];
                
                r_data[299] <= r_data[298];
                
                r_data[300] <= r_data[299];
                
                r_data[301] <= r_data[300];
                
                r_data[302] <= r_data[301];
                
                r_data[303] <= r_data[302];
                
                r_data[304] <= r_data[303];
                
                r_data[305] <= r_data[304];
                
                r_data[306] <= r_data[305];
                
                r_data[307] <= r_data[306];
                
                r_data[308] <= r_data[307];
                
                r_data[309] <= r_data[308];
                
                r_data[310] <= r_data[309];
                
                r_data[311] <= r_data[310];
                
                r_data[312] <= r_data[311];
                
                r_data[313] <= r_data[312];
                
                r_data[314] <= r_data[313];
                
                r_data[315] <= r_data[314];
                
                r_data[316] <= r_data[315];
                
                r_data[317] <= r_data[316];
                
                r_data[318] <= r_data[317];
                
                r_data[319] <= r_data[318];
                
                r_data[320] <= r_data[319];
                
                r_data[321] <= r_data[320];
                
                r_data[322] <= r_data[321];
                
                r_data[323] <= r_data[322];
                
                r_data[324] <= r_data[323];
                
                r_data[325] <= r_data[324];
                
                r_data[326] <= r_data[325];
                
                r_data[327] <= r_data[326];
                
                r_data[328] <= r_data[327];
                
                r_data[329] <= r_data[328];
                
                r_data[330] <= r_data[329];
                
                r_data[331] <= r_data[330];
                
                r_data[332] <= r_data[331];
                
                r_data[333] <= r_data[332];
                
                r_data[334] <= r_data[333];
                
                r_data[335] <= r_data[334];
                
                r_data[336] <= r_data[335];
                
                r_data[337] <= r_data[336];
                
                r_data[338] <= r_data[337];
                
                r_data[339] <= r_data[338];
                
                r_data[340] <= r_data[339];
                
                r_data[341] <= r_data[340];
                
                r_data[342] <= r_data[341];
                
                r_data[343] <= r_data[342];
                
                r_data[344] <= r_data[343];
                
                r_data[345] <= r_data[344];
                
                r_data[346] <= r_data[345];
                
                r_data[347] <= r_data[346];
                
                r_data[348] <= r_data[347];
                
                r_data[349] <= r_data[348];
                
                r_data[350] <= r_data[349];
                
                r_data[351] <= r_data[350];
                
                r_data[352] <= r_data[351];
                
                r_data[353] <= r_data[352];
                
                r_data[354] <= r_data[353];
                
                r_data[355] <= r_data[354];
                
                r_data[356] <= r_data[355];
                
                r_data[357] <= r_data[356];
                
                r_data[358] <= r_data[357];
                
                r_data[359] <= r_data[358];
                
                r_data[360] <= r_data[359];
                
                r_data[361] <= r_data[360];
                
                r_data[362] <= r_data[361];
                
                r_data[363] <= r_data[362];
                
                r_data[364] <= r_data[363];
                
                r_data[365] <= r_data[364];
                
                r_data[366] <= r_data[365];
                
                r_data[367] <= r_data[366];
                
                r_data[368] <= r_data[367];
                
                r_data[369] <= r_data[368];
                
                r_data[370] <= r_data[369];
                
                r_data[371] <= r_data[370];
                
                r_data[372] <= r_data[371];
                
                r_data[373] <= r_data[372];
                
                r_data[374] <= r_data[373];
                
                r_data[375] <= r_data[374];
                
                r_data[376] <= r_data[375];
                
                r_data[377] <= r_data[376];
                
                r_data[378] <= r_data[377];
                
                r_data[379] <= r_data[378];
                
                r_data[380] <= r_data[379];
                
                r_data[381] <= r_data[380];
                
                r_data[382] <= r_data[381];
                
                r_data[383] <= r_data[382];
                
                r_data[384] <= r_data[383];
                
                r_data[385] <= r_data[384];
                
                r_data[386] <= r_data[385];
                
                r_data[387] <= r_data[386];
                
                r_data[388] <= r_data[387];
                
                r_data[389] <= r_data[388];
                
                r_data[390] <= r_data[389];
                
                r_data[391] <= r_data[390];
                
                r_data[392] <= r_data[391];
                
                r_data[393] <= r_data[392];
                
                r_data[394] <= r_data[393];
                
                r_data[395] <= r_data[394];
                
                r_data[396] <= r_data[395];
                
                r_data[397] <= r_data[396];
                
                r_data[398] <= r_data[397];
                
                r_data[399] <= r_data[398];
                
                r_data[400] <= r_data[399];
                
                r_data[401] <= r_data[400];
                
                r_data[402] <= r_data[401];
                
                r_data[403] <= r_data[402];
                
                r_data[404] <= r_data[403];
                
                r_data[405] <= r_data[404];
                
                r_data[406] <= r_data[405];
                
                r_data[407] <= r_data[406];
                
                r_data[408] <= r_data[407];
                
                r_data[409] <= r_data[408];
                
                r_data[410] <= r_data[409];
                
                r_data[411] <= r_data[410];
                
                r_data[412] <= r_data[411];
                
                r_data[413] <= r_data[412];
                
                r_data[414] <= r_data[413];
                
                r_data[415] <= r_data[414];
                
                r_data[416] <= r_data[415];
                
                r_data[417] <= r_data[416];
                
                r_data[418] <= r_data[417];
                
                r_data[419] <= r_data[418];
                
                r_data[420] <= r_data[419];
                
                r_data[421] <= r_data[420];
                
                r_data[422] <= r_data[421];
                
                r_data[423] <= r_data[422];
                
                r_data[424] <= r_data[423];
                
                r_data[425] <= r_data[424];
                
                r_data[426] <= r_data[425];
                
                r_data[427] <= r_data[426];
                
                r_data[428] <= r_data[427];
                
                r_data[429] <= r_data[428];
                
                r_data[430] <= r_data[429];
                
                r_data[431] <= r_data[430];
                
                r_data[432] <= r_data[431];
                
                r_data[433] <= r_data[432];
                
                r_data[434] <= r_data[433];
                
                r_data[435] <= r_data[434];
                
                r_data[436] <= r_data[435];
                
                r_data[437] <= r_data[436];
                
                r_data[438] <= r_data[437];
                
                r_data[439] <= r_data[438];
                
                r_data[440] <= r_data[439];
                
                r_data[441] <= r_data[440];
                
                r_data[442] <= r_data[441];
                
                r_data[443] <= r_data[442];
                
                r_data[444] <= r_data[443];
                
                r_data[445] <= r_data[444];
                
                r_data[446] <= r_data[445];
                
                r_data[447] <= r_data[446];
                
                r_data[448] <= r_data[447];
                
                r_data[449] <= r_data[448];
                
                r_data[450] <= r_data[449];
                
                r_data[451] <= r_data[450];
                
                r_data[452] <= r_data[451];
                
                r_data[453] <= r_data[452];
                
                r_data[454] <= r_data[453];
                
                r_data[455] <= r_data[454];
                
                r_data[456] <= r_data[455];
                
                r_data[457] <= r_data[456];
                
                r_data[458] <= r_data[457];
                
                r_data[459] <= r_data[458];
                
                r_data[460] <= r_data[459];
                
                r_data[461] <= r_data[460];
                
                r_data[462] <= r_data[461];
                
                r_data[463] <= r_data[462];
                
                r_data[464] <= r_data[463];
                
                r_data[465] <= r_data[464];
                
                r_data[466] <= r_data[465];
                
                r_data[467] <= r_data[466];
                
                r_data[468] <= r_data[467];
                
                r_data[469] <= r_data[468];
                
                r_data[470] <= r_data[469];
                
                r_data[471] <= r_data[470];
                
                r_data[472] <= r_data[471];
                
                r_data[473] <= r_data[472];
                
                r_data[474] <= r_data[473];
                
                r_data[475] <= r_data[474];
                
                r_data[476] <= r_data[475];
                
                r_data[477] <= r_data[476];
                
                r_data[478] <= r_data[477];
                
                r_data[479] <= r_data[478];
                
                r_data[480] <= r_data[479];
                
                r_data[481] <= r_data[480];
                
                r_data[482] <= r_data[481];
                
                r_data[483] <= r_data[482];
                
                r_data[484] <= r_data[483];
                
                r_data[485] <= r_data[484];
                
                r_data[486] <= r_data[485];
                
                r_data[487] <= r_data[486];
                
                r_data[488] <= r_data[487];
                
                r_data[489] <= r_data[488];
                
                r_data[490] <= r_data[489];
                
                r_data[491] <= r_data[490];
                
                r_data[492] <= r_data[491];
                
                r_data[493] <= r_data[492];
                
                r_data[494] <= r_data[493];
                
                r_data[495] <= r_data[494];
                
                r_data[496] <= r_data[495];
                
                r_data[497] <= r_data[496];
                
                r_data[498] <= r_data[497];
                
                r_data[499] <= r_data[498];
                
                r_data[500] <= r_data[499];
                
                r_data[501] <= r_data[500];
                
                r_data[502] <= r_data[501];
                
                r_data[503] <= r_data[502];
                
                r_data[504] <= r_data[503];
                
                r_data[505] <= r_data[504];
                
                r_data[506] <= r_data[505];
                
                r_data[507] <= r_data[506];
                
                r_data[508] <= r_data[507];
                
                r_data[509] <= r_data[508];
                
                r_data[510] <= r_data[509];
                
                r_data[511] <= r_data[510];
                
                r_data[512] <= r_data[511];
                
                r_data[513] <= r_data[512];
                
                r_data[514] <= r_data[513];
                
                r_data[515] <= r_data[514];
                
                r_data[516] <= r_data[515];
                
                r_data[517] <= r_data[516];
                
                r_data[518] <= r_data[517];
                
                r_data[519] <= r_data[518];
                
                r_data[520] <= r_data[519];
                
                r_data[521] <= r_data[520];
                
                r_data[522] <= r_data[521];
                
                r_data[523] <= r_data[522];
                
                r_data[524] <= r_data[523];
                
                r_data[525] <= r_data[524];
                
                r_data[526] <= r_data[525];
                
                r_data[527] <= r_data[526];
                
                r_data[528] <= r_data[527];
                
                r_data[529] <= r_data[528];
                
                r_data[530] <= r_data[529];
                
                r_data[531] <= r_data[530];
                
                r_data[532] <= r_data[531];
                
                r_data[533] <= r_data[532];
                
                r_data[534] <= r_data[533];
                
                r_data[535] <= r_data[534];
                
                r_data[536] <= r_data[535];
                
                r_data[537] <= r_data[536];
                
                r_data[538] <= r_data[537];
                
                r_data[539] <= r_data[538];
                
                r_data[540] <= r_data[539];
                
                r_data[541] <= r_data[540];
                
                r_data[542] <= r_data[541];
                
                r_data[543] <= r_data[542];
                
                r_data[544] <= r_data[543];
                
                r_data[545] <= r_data[544];
                
                r_data[546] <= r_data[545];
                
                r_data[547] <= r_data[546];
                
                r_data[548] <= r_data[547];
                
                r_data[549] <= r_data[548];
                
                r_data[550] <= r_data[549];
                
                r_data[551] <= r_data[550];
                
                r_data[552] <= r_data[551];
                
                r_data[553] <= r_data[552];
                
                r_data[554] <= r_data[553];
                
                r_data[555] <= r_data[554];
                
                r_data[556] <= r_data[555];
                
                r_data[557] <= r_data[556];
                
                r_data[558] <= r_data[557];
                
                r_data[559] <= r_data[558];
                
                r_data[560] <= r_data[559];
                
                r_data[561] <= r_data[560];
                
                r_data[562] <= r_data[561];
                
                r_data[563] <= r_data[562];
                
                r_data[564] <= r_data[563];
                
                r_data[565] <= r_data[564];
                
                r_data[566] <= r_data[565];
                
                r_data[567] <= r_data[566];
                
                r_data[568] <= r_data[567];
                
                r_data[569] <= r_data[568];
                
                r_data[570] <= r_data[569];
                
                r_data[571] <= r_data[570];
                
                r_data[572] <= r_data[571];
                
                r_data[573] <= r_data[572];
                
                r_data[574] <= r_data[573];
                
                r_data[575] <= r_data[574];
                
                r_data[576] <= r_data[575];
                
                r_data[577] <= r_data[576];
                
                r_data[578] <= r_data[577];
                
                r_data[579] <= r_data[578];
                
                r_data[580] <= r_data[579];
                
                r_data[581] <= r_data[580];
                
                r_data[582] <= r_data[581];
                
                r_data[583] <= r_data[582];
                
                r_data[584] <= r_data[583];
                
                r_data[585] <= r_data[584];
                
                r_data[586] <= r_data[585];
                
                r_data[587] <= r_data[586];
                
                r_data[588] <= r_data[587];
                
                r_data[589] <= r_data[588];
                
                r_data[590] <= r_data[589];
                
                r_data[591] <= r_data[590];
                
                r_data[592] <= r_data[591];
                
                r_data[593] <= r_data[592];
                
                r_data[594] <= r_data[593];
                
                r_data[595] <= r_data[594];
                
                r_data[596] <= r_data[595];
                
                r_data[597] <= r_data[596];
                
                r_data[598] <= r_data[597];
                
                r_data[599] <= r_data[598];
                
                r_data[600] <= r_data[599];
                
                r_data[601] <= r_data[600];
                
                r_data[602] <= r_data[601];
                
                r_data[603] <= r_data[602];
                
                r_data[604] <= r_data[603];
                
                r_data[605] <= r_data[604];
                
                r_data[606] <= r_data[605];
                
                r_data[607] <= r_data[606];
                
                r_data[608] <= r_data[607];
                
                r_data[609] <= r_data[608];
                
                r_data[610] <= r_data[609];
                
                r_data[611] <= r_data[610];
                
                r_data[612] <= r_data[611];
                
                r_data[613] <= r_data[612];
                
                r_data[614] <= r_data[613];
                
                r_data[615] <= r_data[614];
                
                r_data[616] <= r_data[615];
                
                r_data[617] <= r_data[616];
                
                r_data[618] <= r_data[617];
                
                r_data[619] <= r_data[618];
                
                r_data[620] <= r_data[619];
                
                r_data[621] <= r_data[620];
                
                r_data[622] <= r_data[621];
                
                r_data[623] <= r_data[622];
                
                r_data[624] <= r_data[623];
                
                r_data[625] <= r_data[624];
                
                r_data[626] <= r_data[625];
                
                r_data[627] <= r_data[626];
                
                r_data[628] <= r_data[627];
                
                r_data[629] <= r_data[628];
                
                r_data[630] <= r_data[629];
                
                r_data[631] <= r_data[630];
                
                r_data[632] <= r_data[631];
                
                r_data[633] <= r_data[632];
                
                r_data[634] <= r_data[633];
                
                r_data[635] <= r_data[634];
                
                r_data[636] <= r_data[635];
                
                r_data[637] <= r_data[636];
                
                r_data[638] <= r_data[637];
                
                r_data[639] <= r_data[638];
                
                r_data[640] <= r_data[639];
                
                r_data[641] <= r_data[640];
                
                r_data[642] <= r_data[641];
                
                r_data[643] <= r_data[642];
                
                r_data[644] <= r_data[643];
                
                r_data[645] <= r_data[644];
                
                r_data[646] <= r_data[645];
                
                r_data[647] <= r_data[646];
                
                r_data[648] <= r_data[647];
                
                r_data[649] <= r_data[648];
                
                r_data[650] <= r_data[649];
                
                r_data[651] <= r_data[650];
                
                r_data[652] <= r_data[651];
                
                r_data[653] <= r_data[652];
                
                r_data[654] <= r_data[653];
                
                r_data[655] <= r_data[654];
                
                r_data[656] <= r_data[655];
                
                r_data[657] <= r_data[656];
                
                r_data[658] <= r_data[657];
                
                r_data[659] <= r_data[658];
                
                r_data[660] <= r_data[659];
                
                r_data[661] <= r_data[660];
                
                r_data[662] <= r_data[661];
                
                r_data[663] <= r_data[662];
                
                r_data[664] <= r_data[663];
                
                r_data[665] <= r_data[664];
                
                r_data[666] <= r_data[665];
                
                r_data[667] <= r_data[666];
                
                r_data[668] <= r_data[667];
                
                r_data[669] <= r_data[668];
                
                r_data[670] <= r_data[669];
                
                r_data[671] <= r_data[670];
                
                r_data[672] <= r_data[671];
                
                r_data[673] <= r_data[672];
                
                r_data[674] <= r_data[673];
                
                r_data[675] <= r_data[674];
                
                r_data[676] <= r_data[675];
                
                r_data[677] <= r_data[676];
                
                r_data[678] <= r_data[677];
                
                r_data[679] <= r_data[678];
                
                r_data[680] <= r_data[679];
                
                r_data[681] <= r_data[680];
                
                r_data[682] <= r_data[681];
                
                r_data[683] <= r_data[682];
                
                r_data[684] <= r_data[683];
                
                r_data[685] <= r_data[684];
                
                r_data[686] <= r_data[685];
                
                r_data[687] <= r_data[686];
                
                r_data[688] <= r_data[687];
                
                r_data[689] <= r_data[688];
                
                r_data[690] <= r_data[689];
                
                r_data[691] <= r_data[690];
                
                r_data[692] <= r_data[691];
                
                r_data[693] <= r_data[692];
                
                r_data[694] <= r_data[693];
                
                r_data[695] <= r_data[694];
                
                r_data[696] <= r_data[695];
                
                r_data[697] <= r_data[696];
                
                r_data[698] <= r_data[697];
                
                r_data[699] <= r_data[698];
                
                r_data[700] <= r_data[699];
                
                r_data[701] <= r_data[700];
                
                r_data[702] <= r_data[701];
                
                r_data[703] <= r_data[702];
                
                r_data[704] <= r_data[703];
                
                r_data[705] <= r_data[704];
                
                r_data[706] <= r_data[705];
                
                r_data[707] <= r_data[706];
                
                r_data[708] <= r_data[707];
                
                r_data[709] <= r_data[708];
                
                r_data[710] <= r_data[709];
                
                r_data[711] <= r_data[710];
                
                r_data[712] <= r_data[711];
                
                r_data[713] <= r_data[712];
                
                r_data[714] <= r_data[713];
                
                r_data[715] <= r_data[714];
                
                r_data[716] <= r_data[715];
                
                r_data[717] <= r_data[716];
                
                r_data[718] <= r_data[717];
                
                r_data[719] <= r_data[718];
                
                r_data[720] <= r_data[719];
                
                r_data[721] <= r_data[720];
                
                r_data[722] <= r_data[721];
                
                r_data[723] <= r_data[722];
                
                r_data[724] <= r_data[723];
                
                r_data[725] <= r_data[724];
                
                r_data[726] <= r_data[725];
                
                r_data[727] <= r_data[726];
                
                r_data[728] <= r_data[727];
                
                r_data[729] <= r_data[728];
                
                r_data[730] <= r_data[729];
                
                r_data[731] <= r_data[730];
                
                r_data[732] <= r_data[731];
                
                r_data[733] <= r_data[732];
                
                r_data[734] <= r_data[733];
                
                r_data[735] <= r_data[734];
                
                r_data[736] <= r_data[735];
                
                r_data[737] <= r_data[736];
                
                r_data[738] <= r_data[737];
                
                r_data[739] <= r_data[738];
                
                r_data[740] <= r_data[739];
                
                r_data[741] <= r_data[740];
                
                r_data[742] <= r_data[741];
                
                r_data[743] <= r_data[742];
                
                r_data[744] <= r_data[743];
                
                r_data[745] <= r_data[744];
                
                r_data[746] <= r_data[745];
                
                r_data[747] <= r_data[746];
                
                r_data[748] <= r_data[747];
                
                r_data[749] <= r_data[748];
                
                r_data[750] <= r_data[749];
                
                r_data[751] <= r_data[750];
                
                r_data[752] <= r_data[751];
                
                r_data[753] <= r_data[752];
                
                r_data[754] <= r_data[753];
                
                r_data[755] <= r_data[754];
                
                r_data[756] <= r_data[755];
                
                r_data[757] <= r_data[756];
                
                r_data[758] <= r_data[757];
                
                r_data[759] <= r_data[758];
                
                r_data[760] <= r_data[759];
                
                r_data[761] <= r_data[760];
                
                r_data[762] <= r_data[761];
                
                r_data[763] <= r_data[762];
                
                r_data[764] <= r_data[763];
                
                r_data[765] <= r_data[764];
                
                r_data[766] <= r_data[765];
                
                r_data[767] <= r_data[766];
                
                r_data[768] <= r_data[767];
                
                r_data[769] <= r_data[768];
                
                r_data[770] <= r_data[769];
                
                r_data[771] <= r_data[770];
                
                r_data[772] <= r_data[771];
                
                r_data[773] <= r_data[772];
                
                r_data[774] <= r_data[773];
                
                r_data[775] <= r_data[774];
                
                r_data[776] <= r_data[775];
                
                r_data[777] <= r_data[776];
                
                r_data[778] <= r_data[777];
                
                r_data[779] <= r_data[778];
                
                r_data[780] <= r_data[779];
                
                r_data[781] <= r_data[780];
                
                r_data[782] <= r_data[781];
                
                r_data[783] <= r_data[782];
                
                r_data[784] <= r_data[783];
                
                r_data[785] <= r_data[784];
                
                r_data[786] <= r_data[785];
                
                r_data[787] <= r_data[786];
                
                r_data[788] <= r_data[787];
                
                r_data[789] <= r_data[788];
                
                r_data[790] <= r_data[789];
                
                r_data[791] <= r_data[790];
                
                r_data[792] <= r_data[791];
                
                r_data[793] <= r_data[792];
                
                r_data[794] <= r_data[793];
                
                r_data[795] <= r_data[794];
                
                r_data[796] <= r_data[795];
                
                r_data[797] <= r_data[796];
                
                r_data[798] <= r_data[797];
                
                r_data[799] <= r_data[798];
                
                r_data[800] <= r_data[799];
                
                r_data[801] <= r_data[800];
                
                r_data[802] <= r_data[801];
                
                r_data[803] <= r_data[802];
                
                r_data[804] <= r_data[803];
                
                r_data[805] <= r_data[804];
                
                r_data[806] <= r_data[805];
                
                r_data[807] <= r_data[806];
                
                r_data[808] <= r_data[807];
                
                r_data[809] <= r_data[808];
                
                r_data[810] <= r_data[809];
                
                r_data[811] <= r_data[810];
                
                r_data[812] <= r_data[811];
                
                r_data[813] <= r_data[812];
                
                r_data[814] <= r_data[813];
                
                r_data[815] <= r_data[814];
                
                r_data[816] <= r_data[815];
                
                r_data[817] <= r_data[816];
                
                r_data[818] <= r_data[817];
                
                r_data[819] <= r_data[818];
                
                r_data[820] <= r_data[819];
                
                r_data[821] <= r_data[820];
                
                r_data[822] <= r_data[821];
                
                r_data[823] <= r_data[822];
                
                r_data[824] <= r_data[823];
                
                r_data[825] <= r_data[824];
                
                r_data[826] <= r_data[825];
                
                r_data[827] <= r_data[826];
                
                r_data[828] <= r_data[827];
                
                r_data[829] <= r_data[828];
                
                r_data[830] <= r_data[829];
                
                r_data[831] <= r_data[830];
                
                r_data[832] <= r_data[831];
                
                r_data[833] <= r_data[832];
                
                r_data[834] <= r_data[833];
                
                r_data[835] <= r_data[834];
                
                r_data[836] <= r_data[835];
                
                r_data[837] <= r_data[836];
                
                r_data[838] <= r_data[837];
                
                r_data[839] <= r_data[838];
                
                r_data[840] <= r_data[839];
                
                r_data[841] <= r_data[840];
                
                r_data[842] <= r_data[841];
                
                r_data[843] <= r_data[842];
                
                r_data[844] <= r_data[843];
                
                r_data[845] <= r_data[844];
                
                r_data[846] <= r_data[845];
                
                r_data[847] <= r_data[846];
                
                r_data[848] <= r_data[847];
                
                r_data[849] <= r_data[848];
                
                r_data[850] <= r_data[849];
                
                r_data[851] <= r_data[850];
                
                r_data[852] <= r_data[851];
                
                r_data[853] <= r_data[852];
                
                r_data[854] <= r_data[853];
                
                r_data[855] <= r_data[854];
                
                r_data[856] <= r_data[855];
                
                r_data[857] <= r_data[856];
                
                r_data[858] <= r_data[857];
                
                r_data[859] <= r_data[858];
                
                r_data[860] <= r_data[859];
                
                r_data[861] <= r_data[860];
                
                r_data[862] <= r_data[861];
                
                r_data[863] <= r_data[862];
                
                r_data[864] <= r_data[863];
                
                r_data[865] <= r_data[864];
                
                r_data[866] <= r_data[865];
                
                r_data[867] <= r_data[866];
                
                r_data[868] <= r_data[867];
                
                r_data[869] <= r_data[868];
                
                r_data[870] <= r_data[869];
                
                r_data[871] <= r_data[870];
                
                r_data[872] <= r_data[871];
                
                r_data[873] <= r_data[872];
                
                r_data[874] <= r_data[873];
                
                r_data[875] <= r_data[874];
                
                r_data[876] <= r_data[875];
                
                r_data[877] <= r_data[876];
                
                r_data[878] <= r_data[877];
                
                r_data[879] <= r_data[878];
                
                r_data[880] <= r_data[879];
                
                r_data[881] <= r_data[880];
                
                r_data[882] <= r_data[881];
                
                r_data[883] <= r_data[882];
                
                r_data[884] <= r_data[883];
                
                r_data[885] <= r_data[884];
                
                r_data[886] <= r_data[885];
                
                r_data[887] <= r_data[886];
                
                r_data[888] <= r_data[887];
                
                r_data[889] <= r_data[888];
                
                r_data[890] <= r_data[889];
                
                r_data[891] <= r_data[890];
                
                r_data[892] <= r_data[891];
                
                r_data[893] <= r_data[892];
                
                r_data[894] <= r_data[893];
                
                r_data[895] <= r_data[894];
                
                r_data[896] <= r_data[895];
                
                r_data[897] <= r_data[896];
                
                r_data[898] <= r_data[897];
                
                r_data[899] <= r_data[898];
                
                r_data[900] <= r_data[899];
                
                r_data[901] <= r_data[900];
                
                r_data[902] <= r_data[901];
                
                r_data[903] <= r_data[902];
                
                r_data[904] <= r_data[903];
                
                r_data[905] <= r_data[904];
                
                r_data[906] <= r_data[905];
                
                r_data[907] <= r_data[906];
                
                r_data[908] <= r_data[907];
                
                r_data[909] <= r_data[908];
                
                r_data[910] <= r_data[909];
                
                r_data[911] <= r_data[910];
                
                r_data[912] <= r_data[911];
                
                r_data[913] <= r_data[912];
                
                r_data[914] <= r_data[913];
                
                r_data[915] <= r_data[914];
                
                r_data[916] <= r_data[915];
                
                r_data[917] <= r_data[916];
                
                r_data[918] <= r_data[917];
                
                r_data[919] <= r_data[918];
                
                r_data[920] <= r_data[919];
                
                r_data[921] <= r_data[920];
                
                r_data[922] <= r_data[921];
                
                r_data[923] <= r_data[922];
                
                r_data[924] <= r_data[923];
                
                r_data[925] <= r_data[924];
                
                r_data[926] <= r_data[925];
                
                r_data[927] <= r_data[926];
                
                r_data[928] <= r_data[927];
                
                r_data[929] <= r_data[928];
                
                r_data[930] <= r_data[929];
                
                r_data[931] <= r_data[930];
                
                r_data[932] <= r_data[931];
                
                r_data[933] <= r_data[932];
                
                r_data[934] <= r_data[933];
                
                r_data[935] <= r_data[934];
                
                r_data[936] <= r_data[935];
                
                r_data[937] <= r_data[936];
                
                r_data[938] <= r_data[937];
                
                r_data[939] <= r_data[938];
                
                r_data[940] <= r_data[939];
                
                r_data[941] <= r_data[940];
                
                r_data[942] <= r_data[941];
                
                r_data[943] <= r_data[942];
                
                r_data[944] <= r_data[943];
                
                r_data[945] <= r_data[944];
                
                r_data[946] <= r_data[945];
                
                r_data[947] <= r_data[946];
                
                r_data[948] <= r_data[947];
                
                r_data[949] <= r_data[948];
                
                r_data[950] <= r_data[949];
                
                r_data[951] <= r_data[950];
                
                r_data[952] <= r_data[951];
                
                r_data[953] <= r_data[952];
                
                r_data[954] <= r_data[953];
                
                r_data[955] <= r_data[954];
                
                r_data[956] <= r_data[955];
                
                r_data[957] <= r_data[956];
                
                r_data[958] <= r_data[957];
                
                r_data[959] <= r_data[958];
                
                r_data[960] <= r_data[959];
                
                r_data[961] <= r_data[960];
                
                r_data[962] <= r_data[961];
                
                r_data[963] <= r_data[962];
                
                r_data[964] <= r_data[963];
                
                r_data[965] <= r_data[964];
                
                r_data[966] <= r_data[965];
                
                r_data[967] <= r_data[966];
                
                r_data[968] <= r_data[967];
                
                r_data[969] <= r_data[968];
                
                r_data[970] <= r_data[969];
                
                r_data[971] <= r_data[970];
                
                r_data[972] <= r_data[971];
                
                r_data[973] <= r_data[972];
                
                r_data[974] <= r_data[973];
                
                r_data[975] <= r_data[974];
                
                r_data[976] <= r_data[975];
                
                r_data[977] <= r_data[976];
                
                r_data[978] <= r_data[977];
                
                r_data[979] <= r_data[978];
                
                r_data[980] <= r_data[979];
                
                r_data[981] <= r_data[980];
                
                r_data[982] <= r_data[981];
                
                r_data[983] <= r_data[982];
                
                r_data[984] <= r_data[983];
                
                r_data[985] <= r_data[984];
                
                r_data[986] <= r_data[985];
                
                r_data[987] <= r_data[986];
                
                r_data[988] <= r_data[987];
                
                r_data[989] <= r_data[988];
                
                r_data[990] <= r_data[989];
                
                r_data[991] <= r_data[990];
                
                r_data[992] <= r_data[991];
                
                r_data[993] <= r_data[992];
                
                r_data[994] <= r_data[993];
                
                r_data[995] <= r_data[994];
                
                r_data[996] <= r_data[995];
                
                r_data[997] <= r_data[996];
                
                r_data[998] <= r_data[997];
                
                r_data[999] <= r_data[998];
                
                r_data[1000] <= r_data[999];
                
                r_data[1001] <= r_data[1000];
                
                r_data[1002] <= r_data[1001];
                
                r_data[1003] <= r_data[1002];
                
                r_data[1004] <= r_data[1003];
                
                r_data[1005] <= r_data[1004];
                
                r_data[1006] <= r_data[1005];
                
                r_data[1007] <= r_data[1006];
                
                r_data[1008] <= r_data[1007];
                
                r_data[1009] <= r_data[1008];
                
                r_data[1010] <= r_data[1009];
                
                r_data[1011] <= r_data[1010];
                
                r_data[1012] <= r_data[1011];
                
                r_data[1013] <= r_data[1012];
                
                r_data[1014] <= r_data[1013];
                
                r_data[1015] <= r_data[1014];
                
                r_data[1016] <= r_data[1015];
                
                r_data[1017] <= r_data[1016];
                
                r_data[1018] <= r_data[1017];
                
                r_data[1019] <= r_data[1018];
                
                r_data[1020] <= r_data[1019];
                
                r_data[1021] <= r_data[1020];
                
                r_data[1022] <= r_data[1021];
                
                r_data[1023] <= r_data[1022];
                
                r_data[1024] <= r_data[1023];
                
                r_data[1025] <= r_data[1024];
                
                r_data[1026] <= r_data[1025];
                
                r_data[1027] <= r_data[1026];
                
                r_data[1028] <= r_data[1027];
                
                r_data[1029] <= r_data[1028];
                
                r_data[1030] <= r_data[1029];
                
                r_data[1031] <= r_data[1030];
                
                r_data[1032] <= r_data[1031];
                
                r_data[1033] <= r_data[1032];
                
                r_data[1034] <= r_data[1033];
                
                r_data[1035] <= r_data[1034];
                
                r_data[1036] <= r_data[1035];
                
                r_data[1037] <= r_data[1036];
                
                r_data[1038] <= r_data[1037];
                
                r_data[1039] <= r_data[1038];
                
                r_data[1040] <= r_data[1039];
                
                r_data[1041] <= r_data[1040];
                
                r_data[1042] <= r_data[1041];
                
                r_data[1043] <= r_data[1042];
                
                r_data[1044] <= r_data[1043];
                
                r_data[1045] <= r_data[1044];
                
                r_data[1046] <= r_data[1045];
                
                r_data[1047] <= r_data[1046];
                
                r_data[1048] <= r_data[1047];
                
                r_data[1049] <= r_data[1048];
                
                r_data[1050] <= r_data[1049];
                
                r_data[1051] <= r_data[1050];
                
                r_data[1052] <= r_data[1051];
                
                r_data[1053] <= r_data[1052];
                
                r_data[1054] <= r_data[1053];
                
                r_data[1055] <= r_data[1054];
                
                r_data[1056] <= r_data[1055];
                
                r_data[1057] <= r_data[1056];
                
                r_data[1058] <= r_data[1057];
                
                r_data[1059] <= r_data[1058];
                
                r_data[1060] <= r_data[1059];
                
                r_data[1061] <= r_data[1060];
                
                r_data[1062] <= r_data[1061];
                
                r_data[1063] <= r_data[1062];
                
                r_data[1064] <= r_data[1063];
                
                r_data[1065] <= r_data[1064];
                
                r_data[1066] <= r_data[1065];
                
                r_data[1067] <= r_data[1066];
                
                r_data[1068] <= r_data[1067];
                
                r_data[1069] <= r_data[1068];
                
                r_data[1070] <= r_data[1069];
                
                r_data[1071] <= r_data[1070];
                
                r_data[1072] <= r_data[1071];
                
                r_data[1073] <= r_data[1072];
                
                r_data[1074] <= r_data[1073];
                
                r_data[1075] <= r_data[1074];
                
                r_data[1076] <= r_data[1075];
                
                r_data[1077] <= r_data[1076];
                
                r_data[1078] <= r_data[1077];
                
                r_data[1079] <= r_data[1078];
                
                r_data[1080] <= r_data[1079];
                
                r_data[1081] <= r_data[1080];
                
                r_data[1082] <= r_data[1081];
                
                r_data[1083] <= r_data[1082];
                
                r_data[1084] <= r_data[1083];
                
                r_data[1085] <= r_data[1084];
                
                r_data[1086] <= r_data[1085];
                
                r_data[1087] <= r_data[1086];
                
                r_data[1088] <= r_data[1087];
                
                r_data[1089] <= r_data[1088];
                
                r_data[1090] <= r_data[1089];
                
                r_data[1091] <= r_data[1090];
                
                r_data[1092] <= r_data[1091];
                
                r_data[1093] <= r_data[1092];
                
                r_data[1094] <= r_data[1093];
                
                r_data[1095] <= r_data[1094];
                
                r_data[1096] <= r_data[1095];
                
                r_data[1097] <= r_data[1096];
                
                r_data[1098] <= r_data[1097];
                
                r_data[1099] <= r_data[1098];
                
                r_data[1100] <= r_data[1099];
                
                r_data[1101] <= r_data[1100];
                
                r_data[1102] <= r_data[1101];
                
                r_data[1103] <= r_data[1102];
                
                r_data[1104] <= r_data[1103];
                
                r_data[1105] <= r_data[1104];
                
                r_data[1106] <= r_data[1105];
                
                r_data[1107] <= r_data[1106];
                
                r_data[1108] <= r_data[1107];
                
                r_data[1109] <= r_data[1108];
                
                r_data[1110] <= r_data[1109];
                
                r_data[1111] <= r_data[1110];
                
                r_data[1112] <= r_data[1111];
                
                r_data[1113] <= r_data[1112];
                
                r_data[1114] <= r_data[1113];
                
                r_data[1115] <= r_data[1114];
                
                r_data[1116] <= r_data[1115];
                
                r_data[1117] <= r_data[1116];
                
                r_data[1118] <= r_data[1117];
                
                r_data[1119] <= r_data[1118];
                
                r_data[1120] <= r_data[1119];
                
                r_data[1121] <= r_data[1120];
                
                r_data[1122] <= r_data[1121];
                
                r_data[1123] <= r_data[1122];
                
                r_data[1124] <= r_data[1123];
                
                r_data[1125] <= r_data[1124];
                
                r_data[1126] <= r_data[1125];
                
                r_data[1127] <= r_data[1126];
                
                r_data[1128] <= r_data[1127];
                
                r_data[1129] <= r_data[1128];
                
                r_data[1130] <= r_data[1129];
                
                r_data[1131] <= r_data[1130];
                
                r_data[1132] <= r_data[1131];
                
                r_data[1133] <= r_data[1132];
                
                r_data[1134] <= r_data[1133];
                
                r_data[1135] <= r_data[1134];
                
                r_data[1136] <= r_data[1135];
                
                r_data[1137] <= r_data[1136];
                
                r_data[1138] <= r_data[1137];
                
                r_data[1139] <= r_data[1138];
                
                r_data[1140] <= r_data[1139];
                
                r_data[1141] <= r_data[1140];
                
                r_data[1142] <= r_data[1141];
                
                r_data[1143] <= r_data[1142];
                
                r_data[1144] <= r_data[1143];
                
                r_data[1145] <= r_data[1144];
                
                r_data[1146] <= r_data[1145];
                
                r_data[1147] <= r_data[1146];
                
                r_data[1148] <= r_data[1147];
                
                r_data[1149] <= r_data[1148];
                
                r_data[1150] <= r_data[1149];
                
                r_data[1151] <= r_data[1150];
                
                r_data[1152] <= r_data[1151];
                
                r_data[1153] <= r_data[1152];
                
                r_data[1154] <= r_data[1153];
                
                r_data[1155] <= r_data[1154];
                
                r_data[1156] <= r_data[1155];
                
                r_data[1157] <= r_data[1156];
                
                r_data[1158] <= r_data[1157];
                
                r_data[1159] <= r_data[1158];
                
                r_data[1160] <= r_data[1159];
                
                r_data[1161] <= r_data[1160];
                
                r_data[1162] <= r_data[1161];
                
                r_data[1163] <= r_data[1162];
                
                r_data[1164] <= r_data[1163];
                
                r_data[1165] <= r_data[1164];
                
                r_data[1166] <= r_data[1165];
                
                r_data[1167] <= r_data[1166];
                
                r_data[1168] <= r_data[1167];
                
                r_data[1169] <= r_data[1168];
                
                r_data[1170] <= r_data[1169];
                
                r_data[1171] <= r_data[1170];
                
                r_data[1172] <= r_data[1171];
                
                r_data[1173] <= r_data[1172];
                
                r_data[1174] <= r_data[1173];
                
                r_data[1175] <= r_data[1174];
                
                r_data[1176] <= r_data[1175];
                
                r_data[1177] <= r_data[1176];
                
                r_data[1178] <= r_data[1177];
                
                r_data[1179] <= r_data[1178];
                
                r_data[1180] <= r_data[1179];
                
                r_data[1181] <= r_data[1180];
                
                r_data[1182] <= r_data[1181];
                
                r_data[1183] <= r_data[1182];
                
                r_data[1184] <= r_data[1183];
                
                r_data[1185] <= r_data[1184];
                
                r_data[1186] <= r_data[1185];
                
                r_data[1187] <= r_data[1186];
                
                r_data[1188] <= r_data[1187];
                
                r_data[1189] <= r_data[1188];
                
                r_data[1190] <= r_data[1189];
                
                r_data[1191] <= r_data[1190];
                
                r_data[1192] <= r_data[1191];
                
                r_data[1193] <= r_data[1192];
                
                r_data[1194] <= r_data[1193];
                
                r_data[1195] <= r_data[1194];
                
                r_data[1196] <= r_data[1195];
                
                r_data[1197] <= r_data[1196];
                
                r_data[1198] <= r_data[1197];
                
                r_data[1199] <= r_data[1198];
                
                r_data[1200] <= r_data[1199];
                
                r_data[1201] <= r_data[1200];
                
                r_data[1202] <= r_data[1201];
                
                r_data[1203] <= r_data[1202];
                
                r_data[1204] <= r_data[1203];
                
                r_data[1205] <= r_data[1204];
                
                r_data[1206] <= r_data[1205];
                
                r_data[1207] <= r_data[1206];
                
                r_data[1208] <= r_data[1207];
                
                r_data[1209] <= r_data[1208];
                
                r_data[1210] <= r_data[1209];
                
                r_data[1211] <= r_data[1210];
                
                r_data[1212] <= r_data[1211];
                
                r_data[1213] <= r_data[1212];
                
                r_data[1214] <= r_data[1213];
                
                r_data[1215] <= r_data[1214];
                
                r_data[1216] <= r_data[1215];
                
                r_data[1217] <= r_data[1216];
                
                r_data[1218] <= r_data[1217];
                
                r_data[1219] <= r_data[1218];
                
                r_data[1220] <= r_data[1219];
                
                r_data[1221] <= r_data[1220];
                
                r_data[1222] <= r_data[1221];
                
                r_data[1223] <= r_data[1222];
                
                r_data[1224] <= r_data[1223];
                
                r_data[1225] <= r_data[1224];
                
                r_data[1226] <= r_data[1225];
                
                r_data[1227] <= r_data[1226];
                
                r_data[1228] <= r_data[1227];
                
                r_data[1229] <= r_data[1228];
                
                r_data[1230] <= r_data[1229];
                
                r_data[1231] <= r_data[1230];
                
                r_data[1232] <= r_data[1231];
                
                r_data[1233] <= r_data[1232];
                
                r_data[1234] <= r_data[1233];
                
                r_data[1235] <= r_data[1234];
                
                r_data[1236] <= r_data[1235];
                
                r_data[1237] <= r_data[1236];
                
                r_data[1238] <= r_data[1237];
                
                r_data[1239] <= r_data[1238];
                
                r_data[1240] <= r_data[1239];
                
                r_data[1241] <= r_data[1240];
                
                r_data[1242] <= r_data[1241];
                
                r_data[1243] <= r_data[1242];
                
                r_data[1244] <= r_data[1243];
                
                r_data[1245] <= r_data[1244];
                
                r_data[1246] <= r_data[1245];
                
                r_data[1247] <= r_data[1246];
                
                r_data[1248] <= r_data[1247];
                
                r_data[1249] <= r_data[1248];
                
                r_data[1250] <= r_data[1249];
                
                r_data[1251] <= r_data[1250];
                
                r_data[1252] <= r_data[1251];
                
                r_data[1253] <= r_data[1252];
                
                r_data[1254] <= r_data[1253];
                
                r_data[1255] <= r_data[1254];
                
                r_data[1256] <= r_data[1255];
                
                r_data[1257] <= r_data[1256];
                
                r_data[1258] <= r_data[1257];
                
                r_data[1259] <= r_data[1258];
                
                r_data[1260] <= r_data[1259];
                
                r_data[1261] <= r_data[1260];
                
                r_data[1262] <= r_data[1261];
                
                r_data[1263] <= r_data[1262];
                
                r_data[1264] <= r_data[1263];
                
                r_data[1265] <= r_data[1264];
                
                r_data[1266] <= r_data[1265];
                
                r_data[1267] <= r_data[1266];
                
                r_data[1268] <= r_data[1267];
                
                r_data[1269] <= r_data[1268];
                
                r_data[1270] <= r_data[1269];
                
                r_data[1271] <= r_data[1270];
                
                r_data[1272] <= r_data[1271];
                
                r_data[1273] <= r_data[1272];
                
                r_data[1274] <= r_data[1273];
                
                r_data[1275] <= r_data[1274];
                
                r_data[1276] <= r_data[1275];
                
                r_data[1277] <= r_data[1276];
                
                r_data[1278] <= r_data[1277];
                
                r_data[1279] <= r_data[1278];
                
                r_data[1280] <= r_data[1279];
                
                r_data[1281] <= r_data[1280];
                
                r_data[1282] <= r_data[1281];
                
                r_data[1283] <= r_data[1282];
                
                r_data[1284] <= r_data[1283];
                
                r_data[1285] <= r_data[1284];
                
                r_data[1286] <= r_data[1285];
                
                r_data[1287] <= r_data[1286];
                
                r_data[1288] <= r_data[1287];
                
                r_data[1289] <= r_data[1288];
                
                r_data[1290] <= r_data[1289];
                
                r_data[1291] <= r_data[1290];
                
                r_data[1292] <= r_data[1291];
                
                r_data[1293] <= r_data[1292];
                
                r_data[1294] <= r_data[1293];
                
                r_data[1295] <= r_data[1294];
                
                r_data[1296] <= r_data[1295];
                
                r_data[1297] <= r_data[1296];
                
                r_data[1298] <= r_data[1297];
                
                r_data[1299] <= r_data[1298];
                
                r_data[1300] <= r_data[1299];
                
                r_data[1301] <= r_data[1300];
                
                r_data[1302] <= r_data[1301];
                
                r_data[1303] <= r_data[1302];
                
                r_data[1304] <= r_data[1303];
                
                r_data[1305] <= r_data[1304];
                
                r_data[1306] <= r_data[1305];
                
                r_data[1307] <= r_data[1306];
                
                r_data[1308] <= r_data[1307];
                
                r_data[1309] <= r_data[1308];
                
                r_data[1310] <= r_data[1309];
                
                r_data[1311] <= r_data[1310];
                
                r_data[1312] <= r_data[1311];
                
                r_data[1313] <= r_data[1312];
                
                r_data[1314] <= r_data[1313];
                
                r_data[1315] <= r_data[1314];
                
                r_data[1316] <= r_data[1315];
                
                r_data[1317] <= r_data[1316];
                
                r_data[1318] <= r_data[1317];
                
                r_data[1319] <= r_data[1318];
                
                r_data[1320] <= r_data[1319];
                
                r_data[1321] <= r_data[1320];
                
                r_data[1322] <= r_data[1321];
                
                r_data[1323] <= r_data[1322];
                
                r_data[1324] <= r_data[1323];
                
                r_data[1325] <= r_data[1324];
                
                r_data[1326] <= r_data[1325];
                
                r_data[1327] <= r_data[1326];
                
                r_data[1328] <= r_data[1327];
                
                r_data[1329] <= r_data[1328];
                
                r_data[1330] <= r_data[1329];
                
                r_data[1331] <= r_data[1330];
                
                r_data[1332] <= r_data[1331];
                
                r_data[1333] <= r_data[1332];
                
                r_data[1334] <= r_data[1333];
                
                r_data[1335] <= r_data[1334];
                
                r_data[1336] <= r_data[1335];
                
                r_data[1337] <= r_data[1336];
                
                r_data[1338] <= r_data[1337];
                
                r_data[1339] <= r_data[1338];
                
                r_data[1340] <= r_data[1339];
                
                r_data[1341] <= r_data[1340];
                
                r_data[1342] <= r_data[1341];
                
                r_data[1343] <= r_data[1342];
                
                r_data[1344] <= r_data[1343];
                
                r_data[1345] <= r_data[1344];
                
                r_data[1346] <= r_data[1345];
                
                r_data[1347] <= r_data[1346];
                
                r_data[1348] <= r_data[1347];
                
                r_data[1349] <= r_data[1348];
                
                r_data[1350] <= r_data[1349];
                
                r_data[1351] <= r_data[1350];
                
                r_data[1352] <= r_data[1351];
                
                r_data[1353] <= r_data[1352];
                
                r_data[1354] <= r_data[1353];
                
                r_data[1355] <= r_data[1354];
                
                r_data[1356] <= r_data[1355];
                
                r_data[1357] <= r_data[1356];
                
                r_data[1358] <= r_data[1357];
                
                r_data[1359] <= r_data[1358];
                
                r_data[1360] <= r_data[1359];
                
                r_data[1361] <= r_data[1360];
                
                r_data[1362] <= r_data[1361];
                
                r_data[1363] <= r_data[1362];
                
                r_data[1364] <= r_data[1363];
                
                r_data[1365] <= r_data[1364];
                
                r_data[1366] <= r_data[1365];
                
                r_data[1367] <= r_data[1366];
                
                r_data[1368] <= r_data[1367];
                
                r_data[1369] <= r_data[1368];
                
                r_data[1370] <= r_data[1369];
                
                r_data[1371] <= r_data[1370];
                
                r_data[1372] <= r_data[1371];
                
                r_data[1373] <= r_data[1372];
                
                r_data[1374] <= r_data[1373];
                
                r_data[1375] <= r_data[1374];
                
                r_data[1376] <= r_data[1375];
                
                r_data[1377] <= r_data[1376];
                
                r_data[1378] <= r_data[1377];
                
                r_data[1379] <= r_data[1378];
                
                r_data[1380] <= r_data[1379];
                
                r_data[1381] <= r_data[1380];
                
                r_data[1382] <= r_data[1381];
                
                r_data[1383] <= r_data[1382];
                
                r_data[1384] <= r_data[1383];
                
                r_data[1385] <= r_data[1384];
                
                r_data[1386] <= r_data[1385];
                
                r_data[1387] <= r_data[1386];
                
                r_data[1388] <= r_data[1387];
                
                r_data[1389] <= r_data[1388];
                
                r_data[1390] <= r_data[1389];
                
                r_data[1391] <= r_data[1390];
                
                r_data[1392] <= r_data[1391];
                
                r_data[1393] <= r_data[1392];
                
                r_data[1394] <= r_data[1393];
                
                r_data[1395] <= r_data[1394];
                
                r_data[1396] <= r_data[1395];
                
                r_data[1397] <= r_data[1396];
                
                r_data[1398] <= r_data[1397];
                
                r_data[1399] <= r_data[1398];
                
                r_data[1400] <= r_data[1399];
                
                r_data[1401] <= r_data[1400];
                
                r_data[1402] <= r_data[1401];
                
                r_data[1403] <= r_data[1402];
                
                r_data[1404] <= r_data[1403];
                
                r_data[1405] <= r_data[1404];
                
                r_data[1406] <= r_data[1405];
                
                r_data[1407] <= r_data[1406];
                
                r_data[1408] <= r_data[1407];
                
                r_data[1409] <= r_data[1408];
                
                r_data[1410] <= r_data[1409];
                
                r_data[1411] <= r_data[1410];
                
                r_data[1412] <= r_data[1411];
                
                r_data[1413] <= r_data[1412];
                
                r_data[1414] <= r_data[1413];
                
                r_data[1415] <= r_data[1414];
                
                r_data[1416] <= r_data[1415];
                
                r_data[1417] <= r_data[1416];
                
                r_data[1418] <= r_data[1417];
                
                r_data[1419] <= r_data[1418];
                
                r_data[1420] <= r_data[1419];
                
                r_data[1421] <= r_data[1420];
                
                r_data[1422] <= r_data[1421];
                
                r_data[1423] <= r_data[1422];
                
                r_data[1424] <= r_data[1423];
                
                r_data[1425] <= r_data[1424];
                
                r_data[1426] <= r_data[1425];
                
                r_data[1427] <= r_data[1426];
                
                r_data[1428] <= r_data[1427];
                
                r_data[1429] <= r_data[1428];
                
                r_data[1430] <= r_data[1429];
                
                r_data[1431] <= r_data[1430];
                
                r_data[1432] <= r_data[1431];
                
                r_data[1433] <= r_data[1432];
                
                r_data[1434] <= r_data[1433];
                
                r_data[1435] <= r_data[1434];
                
                r_data[1436] <= r_data[1435];
                
                r_data[1437] <= r_data[1436];
                
                r_data[1438] <= r_data[1437];
                
                r_data[1439] <= r_data[1438];
                
                r_data[1440] <= r_data[1439];
                
                r_data[1441] <= r_data[1440];
                
                r_data[1442] <= r_data[1441];
                
                r_data[1443] <= r_data[1442];
                
                r_data[1444] <= r_data[1443];
                
                r_data[1445] <= r_data[1444];
                
                r_data[1446] <= r_data[1445];
                
                r_data[1447] <= r_data[1446];
                
                r_data[1448] <= r_data[1447];
                
                r_data[1449] <= r_data[1448];
                
                r_data[1450] <= r_data[1449];
                
                r_data[1451] <= r_data[1450];
                
                r_data[1452] <= r_data[1451];
                
                r_data[1453] <= r_data[1452];
                
                r_data[1454] <= r_data[1453];
                
                r_data[1455] <= r_data[1454];
                
                r_data[1456] <= r_data[1455];
                
                r_data[1457] <= r_data[1456];
                
                r_data[1458] <= r_data[1457];
                
                r_data[1459] <= r_data[1458];
                
                r_data[1460] <= r_data[1459];
                
                r_data[1461] <= r_data[1460];
                
                r_data[1462] <= r_data[1461];
                
                r_data[1463] <= r_data[1462];
                
                r_data[1464] <= r_data[1463];
                
                r_data[1465] <= r_data[1464];
                
                r_data[1466] <= r_data[1465];
                
                r_data[1467] <= r_data[1466];
                
                r_data[1468] <= r_data[1467];
                
                r_data[1469] <= r_data[1468];
                
                r_data[1470] <= r_data[1469];
                
                r_data[1471] <= r_data[1470];
                
                r_data[1472] <= r_data[1471];
                
                r_data[1473] <= r_data[1472];
                
                r_data[1474] <= r_data[1473];
                
                r_data[1475] <= r_data[1474];
                
                r_data[1476] <= r_data[1475];
                
                r_data[1477] <= r_data[1476];
                
                r_data[1478] <= r_data[1477];
                
                r_data[1479] <= r_data[1478];
                
                r_data[1480] <= r_data[1479];
                
                r_data[1481] <= r_data[1480];
                
                r_data[1482] <= r_data[1481];
                
                r_data[1483] <= r_data[1482];
                
                r_data[1484] <= r_data[1483];
                
                r_data[1485] <= r_data[1484];
                
                r_data[1486] <= r_data[1485];
                
                r_data[1487] <= r_data[1486];
                
                r_data[1488] <= r_data[1487];
                
                r_data[1489] <= r_data[1488];
                
                r_data[1490] <= r_data[1489];
                
                r_data[1491] <= r_data[1490];
                
                r_data[1492] <= r_data[1491];
                
                r_data[1493] <= r_data[1492];
                
                r_data[1494] <= r_data[1493];
                
                r_data[1495] <= r_data[1494];
                
                r_data[1496] <= r_data[1495];
                
                r_data[1497] <= r_data[1496];
                
                r_data[1498] <= r_data[1497];
                
                r_data[1499] <= r_data[1498];
                
                r_data[1500] <= r_data[1499];
                
                r_data[1501] <= r_data[1500];
                
                r_data[1502] <= r_data[1501];
                
                r_data[1503] <= r_data[1502];
                
                r_data[1504] <= r_data[1503];
                
                r_data[1505] <= r_data[1504];
                
                r_data[1506] <= r_data[1505];
                
                r_data[1507] <= r_data[1506];
                
                r_data[1508] <= r_data[1507];
                
                r_data[1509] <= r_data[1508];
                
                r_data[1510] <= r_data[1509];
                
                r_data[1511] <= r_data[1510];
                
                r_data[1512] <= r_data[1511];
                
                r_data[1513] <= r_data[1512];
                
                r_data[1514] <= r_data[1513];
                
                r_data[1515] <= r_data[1514];
                
                r_data[1516] <= r_data[1515];
                
                r_data[1517] <= r_data[1516];
                
                r_data[1518] <= r_data[1517];
                
                r_data[1519] <= r_data[1518];
                
                r_data[1520] <= r_data[1519];
                
                r_data[1521] <= r_data[1520];
                
                r_data[1522] <= r_data[1521];
                
                r_data[1523] <= r_data[1522];
                
                r_data[1524] <= r_data[1523];
                
                r_data[1525] <= r_data[1524];
                
                r_data[1526] <= r_data[1525];
                
                r_data[1527] <= r_data[1526];
                
                r_data[1528] <= r_data[1527];
                
                r_data[1529] <= r_data[1528];
                
                r_data[1530] <= r_data[1529];
                
                r_data[1531] <= r_data[1530];
                
                r_data[1532] <= r_data[1531];
                
                r_data[1533] <= r_data[1532];
                
                r_data[1534] <= r_data[1533];
                
                r_data[1535] <= r_data[1534];
                
                r_data[1536] <= r_data[1535];
                
                r_data[1537] <= r_data[1536];
                
                r_data[1538] <= r_data[1537];
                
                r_data[1539] <= r_data[1538];
                
                r_data[1540] <= r_data[1539];
                
                r_data[1541] <= r_data[1540];
                
                r_data[1542] <= r_data[1541];
                
                r_data[1543] <= r_data[1542];
                
                r_data[1544] <= r_data[1543];
                
                r_data[1545] <= r_data[1544];
                
                r_data[1546] <= r_data[1545];
                
                r_data[1547] <= r_data[1546];
                
                r_data[1548] <= r_data[1547];
                
                r_data[1549] <= r_data[1548];
                
                r_data[1550] <= r_data[1549];
                
                r_data[1551] <= r_data[1550];
                
                r_data[1552] <= r_data[1551];
                
                r_data[1553] <= r_data[1552];
                
                r_data[1554] <= r_data[1553];
                
                r_data[1555] <= r_data[1554];
                
                r_data[1556] <= r_data[1555];
                
                r_data[1557] <= r_data[1556];
                
                r_data[1558] <= r_data[1557];
                
                r_data[1559] <= r_data[1558];
                
                r_data[1560] <= r_data[1559];
                
                r_data[1561] <= r_data[1560];
                
                r_data[1562] <= r_data[1561];
                
                r_data[1563] <= r_data[1562];
                
                r_data[1564] <= r_data[1563];
                
                r_data[1565] <= r_data[1564];
                
                r_data[1566] <= r_data[1565];
                
                r_data[1567] <= r_data[1566];
                
                r_data[1568] <= r_data[1567];
                
                r_data[1569] <= r_data[1568];
                
                r_data[1570] <= r_data[1569];
                
                r_data[1571] <= r_data[1570];
                
                r_data[1572] <= r_data[1571];
                
                r_data[1573] <= r_data[1572];
                
                r_data[1574] <= r_data[1573];
                
                r_data[1575] <= r_data[1574];
                
                r_data[1576] <= r_data[1575];
                
                r_data[1577] <= r_data[1576];
                
                r_data[1578] <= r_data[1577];
                
                r_data[1579] <= r_data[1578];
                
                r_data[1580] <= r_data[1579];
                
                r_data[1581] <= r_data[1580];
                
                r_data[1582] <= r_data[1581];
                
                r_data[1583] <= r_data[1582];
                
                r_data[1584] <= r_data[1583];
                
                r_data[1585] <= r_data[1584];
                
                r_data[1586] <= r_data[1585];
                
                r_data[1587] <= r_data[1586];
                
                r_data[1588] <= r_data[1587];
                
                r_data[1589] <= r_data[1588];
                
                r_data[1590] <= r_data[1589];
                
                r_data[1591] <= r_data[1590];
                
                r_data[1592] <= r_data[1591];
                
                r_data[1593] <= r_data[1592];
                
                r_data[1594] <= r_data[1593];
                
                r_data[1595] <= r_data[1594];
                
                r_data[1596] <= r_data[1595];
                
                r_data[1597] <= r_data[1596];
                
                r_data[1598] <= r_data[1597];
                
                r_data[1599] <= r_data[1598];
                
                r_data[1600] <= r_data[1599];
                
                r_data[1601] <= r_data[1600];
                
                r_data[1602] <= r_data[1601];
                
                r_data[1603] <= r_data[1602];
                
                r_data[1604] <= r_data[1603];
                
                r_data[1605] <= r_data[1604];
                
                r_data[1606] <= r_data[1605];
                
                r_data[1607] <= r_data[1606];
                
                r_data[1608] <= r_data[1607];
                
                r_data[1609] <= r_data[1608];
                
                r_data[1610] <= r_data[1609];
                
                r_data[1611] <= r_data[1610];
                
                r_data[1612] <= r_data[1611];
                
                r_data[1613] <= r_data[1612];
                
                r_data[1614] <= r_data[1613];
                
                r_data[1615] <= r_data[1614];
                
                r_data[1616] <= r_data[1615];
                
                r_data[1617] <= r_data[1616];
                
                r_data[1618] <= r_data[1617];
                
                r_data[1619] <= r_data[1618];
                
                r_data[1620] <= r_data[1619];
                
                r_data[1621] <= r_data[1620];
                
                r_data[1622] <= r_data[1621];
                
                r_data[1623] <= r_data[1622];
                
                r_data[1624] <= r_data[1623];
                
                r_data[1625] <= r_data[1624];
                
                r_data[1626] <= r_data[1625];
                
                r_data[1627] <= r_data[1626];
                
                r_data[1628] <= r_data[1627];
                
                r_data[1629] <= r_data[1628];
                
                r_data[1630] <= r_data[1629];
                
                r_data[1631] <= r_data[1630];
                
                r_data[1632] <= r_data[1631];
                
                r_data[1633] <= r_data[1632];
                
                r_data[1634] <= r_data[1633];
                
                r_data[1635] <= r_data[1634];
                
                r_data[1636] <= r_data[1635];
                
                r_data[1637] <= r_data[1636];
                
                r_data[1638] <= r_data[1637];
                
                r_data[1639] <= r_data[1638];
                
                r_data[1640] <= r_data[1639];
                
                r_data[1641] <= r_data[1640];
                
                r_data[1642] <= r_data[1641];
                
                r_data[1643] <= r_data[1642];
                
                r_data[1644] <= r_data[1643];
                
                r_data[1645] <= r_data[1644];
                
                r_data[1646] <= r_data[1645];
                
                r_data[1647] <= r_data[1646];
                
                r_data[1648] <= r_data[1647];
                
                r_data[1649] <= r_data[1648];
                
                r_data[1650] <= r_data[1649];
                
                r_data[1651] <= r_data[1650];
                
                r_data[1652] <= r_data[1651];
                
                r_data[1653] <= r_data[1652];
                
                r_data[1654] <= r_data[1653];
                
                r_data[1655] <= r_data[1654];
                
                r_data[1656] <= r_data[1655];
                
                r_data[1657] <= r_data[1656];
                
                r_data[1658] <= r_data[1657];
                
                r_data[1659] <= r_data[1658];
                
                r_data[1660] <= r_data[1659];
                
                r_data[1661] <= r_data[1660];
                
                r_data[1662] <= r_data[1661];
                
                r_data[1663] <= r_data[1662];
                
                r_data[1664] <= r_data[1663];
                
                r_data[1665] <= r_data[1664];
                
                r_data[1666] <= r_data[1665];
                
                r_data[1667] <= r_data[1666];
                
                r_data[1668] <= r_data[1667];
                
                r_data[1669] <= r_data[1668];
                
                r_data[1670] <= r_data[1669];
                
                r_data[1671] <= r_data[1670];
                
                r_data[1672] <= r_data[1671];
                
                r_data[1673] <= r_data[1672];
                
                r_data[1674] <= r_data[1673];
                
                r_data[1675] <= r_data[1674];
                
                r_data[1676] <= r_data[1675];
                
                r_data[1677] <= r_data[1676];
                
                r_data[1678] <= r_data[1677];
                
                r_data[1679] <= r_data[1678];
                
                r_data[1680] <= r_data[1679];
                
                r_data[1681] <= r_data[1680];
                
                r_data[1682] <= r_data[1681];
                
                r_data[1683] <= r_data[1682];
                
                r_data[1684] <= r_data[1683];
                
                r_data[1685] <= r_data[1684];
                
                r_data[1686] <= r_data[1685];
                
                r_data[1687] <= r_data[1686];
                
                r_data[1688] <= r_data[1687];
                
                r_data[1689] <= r_data[1688];
                
                r_data[1690] <= r_data[1689];
                
                r_data[1691] <= r_data[1690];
                
                r_data[1692] <= r_data[1691];
                
                r_data[1693] <= r_data[1692];
                
                r_data[1694] <= r_data[1693];
                
                r_data[1695] <= r_data[1694];
                
                r_data[1696] <= r_data[1695];
                
                r_data[1697] <= r_data[1696];
                
                r_data[1698] <= r_data[1697];
                
                r_data[1699] <= r_data[1698];
                
                r_data[1700] <= r_data[1699];
                
                r_data[1701] <= r_data[1700];
                
                r_data[1702] <= r_data[1701];
                
                r_data[1703] <= r_data[1702];
                
                r_data[1704] <= r_data[1703];
                
                r_data[1705] <= r_data[1704];
                
                r_data[1706] <= r_data[1705];
                
                r_data[1707] <= r_data[1706];
                
                r_data[1708] <= r_data[1707];
                
                r_data[1709] <= r_data[1708];
                
                r_data[1710] <= r_data[1709];
                
                r_data[1711] <= r_data[1710];
                
                r_data[1712] <= r_data[1711];
                
                r_data[1713] <= r_data[1712];
                
                r_data[1714] <= r_data[1713];
                
                r_data[1715] <= r_data[1714];
                
                r_data[1716] <= r_data[1715];
                
                r_data[1717] <= r_data[1716];
                
                r_data[1718] <= r_data[1717];
                
                r_data[1719] <= r_data[1718];
                
                r_data[1720] <= r_data[1719];
                
                r_data[1721] <= r_data[1720];
                
                r_data[1722] <= r_data[1721];
                
                r_data[1723] <= r_data[1722];
                
                r_data[1724] <= r_data[1723];
                
                r_data[1725] <= r_data[1724];
                
                r_data[1726] <= r_data[1725];
                
                r_data[1727] <= r_data[1726];
                
                r_data[1728] <= r_data[1727];
                
                r_data[1729] <= r_data[1728];
                
                r_data[1730] <= r_data[1729];
                
                r_data[1731] <= r_data[1730];
                
                r_data[1732] <= r_data[1731];
                
                r_data[1733] <= r_data[1732];
                
                r_data[1734] <= r_data[1733];
                
                r_data[1735] <= r_data[1734];
                
                r_data[1736] <= r_data[1735];
                
                r_data[1737] <= r_data[1736];
                
                r_data[1738] <= r_data[1737];
                
                r_data[1739] <= r_data[1738];
                
                r_data[1740] <= r_data[1739];
                
                r_data[1741] <= r_data[1740];
                
                r_data[1742] <= r_data[1741];
                
                r_data[1743] <= r_data[1742];
                
                r_data[1744] <= r_data[1743];
                
                r_data[1745] <= r_data[1744];
                
                r_data[1746] <= r_data[1745];
                
                r_data[1747] <= r_data[1746];
                
                r_data[1748] <= r_data[1747];
                
                r_data[1749] <= r_data[1748];
                
                r_data[1750] <= r_data[1749];
                
                r_data[1751] <= r_data[1750];
                
                r_data[1752] <= r_data[1751];
                
                r_data[1753] <= r_data[1752];
                
                r_data[1754] <= r_data[1753];
                
                r_data[1755] <= r_data[1754];
                
                r_data[1756] <= r_data[1755];
                
                r_data[1757] <= r_data[1756];
                
                r_data[1758] <= r_data[1757];
                
                r_data[1759] <= r_data[1758];
                
                r_data[1760] <= r_data[1759];
                
                r_data[1761] <= r_data[1760];
                
                r_data[1762] <= r_data[1761];
                
                r_data[1763] <= r_data[1762];
                
                r_data[1764] <= r_data[1763];
                
                r_data[1765] <= r_data[1764];
                
                r_data[1766] <= r_data[1765];
                
                r_data[1767] <= r_data[1766];
                
                r_data[1768] <= r_data[1767];
                
                r_data[1769] <= r_data[1768];
                
                r_data[1770] <= r_data[1769];
                
                r_data[1771] <= r_data[1770];
                
                r_data[1772] <= r_data[1771];
                
                r_data[1773] <= r_data[1772];
                
                r_data[1774] <= r_data[1773];
                
                r_data[1775] <= r_data[1774];
                
                r_data[1776] <= r_data[1775];
                
                r_data[1777] <= r_data[1776];
                
                r_data[1778] <= r_data[1777];
                
                r_data[1779] <= r_data[1778];
                
                r_data[1780] <= r_data[1779];
                
                r_data[1781] <= r_data[1780];
                
                r_data[1782] <= r_data[1781];
                
                r_data[1783] <= r_data[1782];
                
                r_data[1784] <= r_data[1783];
                
                r_data[1785] <= r_data[1784];
                
                r_data[1786] <= r_data[1785];
                
                r_data[1787] <= r_data[1786];
                
                r_data[1788] <= r_data[1787];
                
                r_data[1789] <= r_data[1788];
                
                r_data[1790] <= r_data[1789];
                
                r_data[1791] <= r_data[1790];
                
                r_data[1792] <= r_data[1791];
                
                r_data[1793] <= r_data[1792];
                
                r_data[1794] <= r_data[1793];
                
                r_data[1795] <= r_data[1794];
                
                r_data[1796] <= r_data[1795];
                
                r_data[1797] <= r_data[1796];
                
                r_data[1798] <= r_data[1797];
                
                r_data[1799] <= r_data[1798];
                
                r_data[1800] <= r_data[1799];
                
                r_data[1801] <= r_data[1800];
                
                r_data[1802] <= r_data[1801];
                
                r_data[1803] <= r_data[1802];
                
                r_data[1804] <= r_data[1803];
                
                r_data[1805] <= r_data[1804];
                
                r_data[1806] <= r_data[1805];
                
                r_data[1807] <= r_data[1806];
                
                r_data[1808] <= r_data[1807];
                
                r_data[1809] <= r_data[1808];
                
                r_data[1810] <= r_data[1809];
                
                r_data[1811] <= r_data[1810];
                
                r_data[1812] <= r_data[1811];
                
                r_data[1813] <= r_data[1812];
                
                r_data[1814] <= r_data[1813];
                
                r_data[1815] <= r_data[1814];
                
                r_data[1816] <= r_data[1815];
                
                r_data[1817] <= r_data[1816];
                
                r_data[1818] <= r_data[1817];
                
                r_data[1819] <= r_data[1818];
                
                r_data[1820] <= r_data[1819];
                
                r_data[1821] <= r_data[1820];
                
                r_data[1822] <= r_data[1821];
                
                r_data[1823] <= r_data[1822];
                
                r_data[1824] <= r_data[1823];
                
                r_data[1825] <= r_data[1824];
                
                r_data[1826] <= r_data[1825];
                
                r_data[1827] <= r_data[1826];
                
                r_data[1828] <= r_data[1827];
                
                r_data[1829] <= r_data[1828];
                
                r_data[1830] <= r_data[1829];
                
                r_data[1831] <= r_data[1830];
                
                r_data[1832] <= r_data[1831];
                
                r_data[1833] <= r_data[1832];
                
                r_data[1834] <= r_data[1833];
                
                r_data[1835] <= r_data[1834];
                
                r_data[1836] <= r_data[1835];
                
                r_data[1837] <= r_data[1836];
                
                r_data[1838] <= r_data[1837];
                
                r_data[1839] <= r_data[1838];
                
                r_data[1840] <= r_data[1839];
                
                r_data[1841] <= r_data[1840];
                
                r_data[1842] <= r_data[1841];
                
                r_data[1843] <= r_data[1842];
                
                r_data[1844] <= r_data[1843];
                
                r_data[1845] <= r_data[1844];
                
                r_data[1846] <= r_data[1845];
                
                r_data[1847] <= r_data[1846];
                
                r_data[1848] <= r_data[1847];
                
                r_data[1849] <= r_data[1848];
                
                r_data[1850] <= r_data[1849];
                
                r_data[1851] <= r_data[1850];
                
                r_data[1852] <= r_data[1851];
                
                r_data[1853] <= r_data[1852];
                
                r_data[1854] <= r_data[1853];
                
                r_data[1855] <= r_data[1854];
                
                r_data[1856] <= r_data[1855];
                
                r_data[1857] <= r_data[1856];
                
                r_data[1858] <= r_data[1857];
                
                r_data[1859] <= r_data[1858];
                
                r_data[1860] <= r_data[1859];
                
                r_data[1861] <= r_data[1860];
                
                r_data[1862] <= r_data[1861];
                
                r_data[1863] <= r_data[1862];
                
                r_data[1864] <= r_data[1863];
                
                r_data[1865] <= r_data[1864];
                
                r_data[1866] <= r_data[1865];
                
                r_data[1867] <= r_data[1866];
                
                r_data[1868] <= r_data[1867];
                
                r_data[1869] <= r_data[1868];
                
                r_data[1870] <= r_data[1869];
                
                r_data[1871] <= r_data[1870];
                
                r_data[1872] <= r_data[1871];
                
                r_data[1873] <= r_data[1872];
                
                r_data[1874] <= r_data[1873];
                
                r_data[1875] <= r_data[1874];
                
                r_data[1876] <= r_data[1875];
                
                r_data[1877] <= r_data[1876];
                
                r_data[1878] <= r_data[1877];
                
                r_data[1879] <= r_data[1878];
                
                r_data[1880] <= r_data[1879];
                
                r_data[1881] <= r_data[1880];
                
                r_data[1882] <= r_data[1881];
                
                r_data[1883] <= r_data[1882];
                
                r_data[1884] <= r_data[1883];
                
                r_data[1885] <= r_data[1884];
                
                r_data[1886] <= r_data[1885];
                
                r_data[1887] <= r_data[1886];
                
                r_data[1888] <= r_data[1887];
                
                r_data[1889] <= r_data[1888];
                
                r_data[1890] <= r_data[1889];
                
                r_data[1891] <= r_data[1890];
                
                r_data[1892] <= r_data[1891];
                
                r_data[1893] <= r_data[1892];
                
                r_data[1894] <= r_data[1893];
                
                r_data[1895] <= r_data[1894];
                
                r_data[1896] <= r_data[1895];
                
                r_data[1897] <= r_data[1896];
                
                r_data[1898] <= r_data[1897];
                
                r_data[1899] <= r_data[1898];
                
                r_data[1900] <= r_data[1899];
                
                r_data[1901] <= r_data[1900];
                
                r_data[1902] <= r_data[1901];
                
                r_data[1903] <= r_data[1902];
                
                r_data[1904] <= r_data[1903];
                
                r_data[1905] <= r_data[1904];
                
                r_data[1906] <= r_data[1905];
                
                r_data[1907] <= r_data[1906];
                
                r_data[1908] <= r_data[1907];
                
                r_data[1909] <= r_data[1908];
                
                r_data[1910] <= r_data[1909];
                
                r_data[1911] <= r_data[1910];
                
                r_data[1912] <= r_data[1911];
                
                r_data[1913] <= r_data[1912];
                
                r_data[1914] <= r_data[1913];
                
                r_data[1915] <= r_data[1914];
                
                r_data[1916] <= r_data[1915];
                
                r_data[1917] <= r_data[1916];
                
                r_data[1918] <= r_data[1917];
                
                r_data[1919] <= r_data[1918];
                
                r_data[1920] <= r_data[1919];
                
                r_data[1921] <= r_data[1920];
                
                r_data[1922] <= r_data[1921];
                
                r_data[1923] <= r_data[1922];
                
                r_data[1924] <= r_data[1923];
                
                r_data[1925] <= r_data[1924];
                
                r_data[1926] <= r_data[1925];
                
                r_data[1927] <= r_data[1926];
                
                r_data[1928] <= r_data[1927];
                
                r_data[1929] <= r_data[1928];
                
                r_data[1930] <= r_data[1929];
                
                r_data[1931] <= r_data[1930];
                
                r_data[1932] <= r_data[1931];
                
                r_data[1933] <= r_data[1932];
                
                r_data[1934] <= r_data[1933];
                
                r_data[1935] <= r_data[1934];
                
                r_data[1936] <= r_data[1935];
                
                r_data[1937] <= r_data[1936];
                
                r_data[1938] <= r_data[1937];
                
                r_data[1939] <= r_data[1938];
                
                r_data[1940] <= r_data[1939];
                
                r_data[1941] <= r_data[1940];
                
                r_data[1942] <= r_data[1941];
                
                r_data[1943] <= r_data[1942];
                
                r_data[1944] <= r_data[1943];
                
                r_data[1945] <= r_data[1944];
                
                r_data[1946] <= r_data[1945];
                
                r_data[1947] <= r_data[1946];
                
                r_data[1948] <= r_data[1947];
                
                r_data[1949] <= r_data[1948];
                
                r_data[1950] <= r_data[1949];
                
                r_data[1951] <= r_data[1950];
                
                r_data[1952] <= r_data[1951];
                
                r_data[1953] <= r_data[1952];
                
                r_data[1954] <= r_data[1953];
                
                r_data[1955] <= r_data[1954];
                
                r_data[1956] <= r_data[1955];
                
                r_data[1957] <= r_data[1956];
                
                r_data[1958] <= r_data[1957];
                
                r_data[1959] <= r_data[1958];
                
                r_data[1960] <= r_data[1959];
                
                r_data[1961] <= r_data[1960];
                
                r_data[1962] <= r_data[1961];
                
                r_data[1963] <= r_data[1962];
                
                r_data[1964] <= r_data[1963];
                
                r_data[1965] <= r_data[1964];
                
                r_data[1966] <= r_data[1965];
                
                r_data[1967] <= r_data[1966];
                
                r_data[1968] <= r_data[1967];
                
                r_data[1969] <= r_data[1968];
                
                r_data[1970] <= r_data[1969];
                
                r_data[1971] <= r_data[1970];
                
                r_data[1972] <= r_data[1971];
                
                r_data[1973] <= r_data[1972];
                
                r_data[1974] <= r_data[1973];
                
                r_data[1975] <= r_data[1974];
                
                r_data[1976] <= r_data[1975];
                
                r_data[1977] <= r_data[1976];
                
                r_data[1978] <= r_data[1977];
                
                r_data[1979] <= r_data[1978];
                
                r_data[1980] <= r_data[1979];
                
                r_data[1981] <= r_data[1980];
                
                r_data[1982] <= r_data[1981];
                
                r_data[1983] <= r_data[1982];
                
                r_data[1984] <= r_data[1983];
                
                r_data[1985] <= r_data[1984];
                
                r_data[1986] <= r_data[1985];
                
                r_data[1987] <= r_data[1986];
                
                r_data[1988] <= r_data[1987];
                
                r_data[1989] <= r_data[1988];
                
                r_data[1990] <= r_data[1989];
                
                r_data[1991] <= r_data[1990];
                
                r_data[1992] <= r_data[1991];
                
                r_data[1993] <= r_data[1992];
                
                r_data[1994] <= r_data[1993];
                
                r_data[1995] <= r_data[1994];
                
                r_data[1996] <= r_data[1995];
                
                r_data[1997] <= r_data[1996];
                
                r_data[1998] <= r_data[1997];
                
                r_data[1999] <= r_data[1998];
                
                r_data[2000] <= r_data[1999];
                
                r_data[2001] <= r_data[2000];
                
                r_data[2002] <= r_data[2001];
                
                r_data[2003] <= r_data[2002];
                
                r_data[2004] <= r_data[2003];
                
                r_data[2005] <= r_data[2004];
                
                r_data[2006] <= r_data[2005];
                
                r_data[2007] <= r_data[2006];
                
                r_data[2008] <= r_data[2007];
                
                r_data[2009] <= r_data[2008];
                
                r_data[2010] <= r_data[2009];
                
                r_data[2011] <= r_data[2010];
                
                r_data[2012] <= r_data[2011];
                
                r_data[2013] <= r_data[2012];
                
                r_data[2014] <= r_data[2013];
                
                r_data[2015] <= r_data[2014];
                
                r_data[2016] <= r_data[2015];
                
                r_data[2017] <= r_data[2016];
                
                r_data[2018] <= r_data[2017];
                
                r_data[2019] <= r_data[2018];
                
                r_data[2020] <= r_data[2019];
                
                r_data[2021] <= r_data[2020];
                
                r_data[2022] <= r_data[2021];
                
                r_data[2023] <= r_data[2022];
                
                r_data[2024] <= r_data[2023];
                
                r_data[2025] <= r_data[2024];
                
                r_data[2026] <= r_data[2025];
                
                r_data[2027] <= r_data[2026];
                
                r_data[2028] <= r_data[2027];
                
                r_data[2029] <= r_data[2028];
                
                r_data[2030] <= r_data[2029];
                
                r_data[2031] <= r_data[2030];
                
                r_data[2032] <= r_data[2031];
                
                r_data[2033] <= r_data[2032];
                
            end
        end
    end
    assign data_out = r_data;   

endmodule