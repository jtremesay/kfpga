module ConfigShiftRegister(
    input data_in,
    output [42367:0] data_out,
    input clock,
    input enable,
    input nreset
);
    reg [42367:0] r_data;
    always @(posedge clock) begin
        if (!nreset) begin
            r_data <= 0;
        end else begin
            if (enable) begin
                
                r_data[0] <= data_in;
                
                r_data[1] <= r_data[0];
                
                r_data[2] <= r_data[1];
                
                r_data[3] <= r_data[2];
                
                r_data[4] <= r_data[3];
                
                r_data[5] <= r_data[4];
                
                r_data[6] <= r_data[5];
                
                r_data[7] <= r_data[6];
                
                r_data[8] <= r_data[7];
                
                r_data[9] <= r_data[8];
                
                r_data[10] <= r_data[9];
                
                r_data[11] <= r_data[10];
                
                r_data[12] <= r_data[11];
                
                r_data[13] <= r_data[12];
                
                r_data[14] <= r_data[13];
                
                r_data[15] <= r_data[14];
                
                r_data[16] <= r_data[15];
                
                r_data[17] <= r_data[16];
                
                r_data[18] <= r_data[17];
                
                r_data[19] <= r_data[18];
                
                r_data[20] <= r_data[19];
                
                r_data[21] <= r_data[20];
                
                r_data[22] <= r_data[21];
                
                r_data[23] <= r_data[22];
                
                r_data[24] <= r_data[23];
                
                r_data[25] <= r_data[24];
                
                r_data[26] <= r_data[25];
                
                r_data[27] <= r_data[26];
                
                r_data[28] <= r_data[27];
                
                r_data[29] <= r_data[28];
                
                r_data[30] <= r_data[29];
                
                r_data[31] <= r_data[30];
                
                r_data[32] <= r_data[31];
                
                r_data[33] <= r_data[32];
                
                r_data[34] <= r_data[33];
                
                r_data[35] <= r_data[34];
                
                r_data[36] <= r_data[35];
                
                r_data[37] <= r_data[36];
                
                r_data[38] <= r_data[37];
                
                r_data[39] <= r_data[38];
                
                r_data[40] <= r_data[39];
                
                r_data[41] <= r_data[40];
                
                r_data[42] <= r_data[41];
                
                r_data[43] <= r_data[42];
                
                r_data[44] <= r_data[43];
                
                r_data[45] <= r_data[44];
                
                r_data[46] <= r_data[45];
                
                r_data[47] <= r_data[46];
                
                r_data[48] <= r_data[47];
                
                r_data[49] <= r_data[48];
                
                r_data[50] <= r_data[49];
                
                r_data[51] <= r_data[50];
                
                r_data[52] <= r_data[51];
                
                r_data[53] <= r_data[52];
                
                r_data[54] <= r_data[53];
                
                r_data[55] <= r_data[54];
                
                r_data[56] <= r_data[55];
                
                r_data[57] <= r_data[56];
                
                r_data[58] <= r_data[57];
                
                r_data[59] <= r_data[58];
                
                r_data[60] <= r_data[59];
                
                r_data[61] <= r_data[60];
                
                r_data[62] <= r_data[61];
                
                r_data[63] <= r_data[62];
                
                r_data[64] <= r_data[63];
                
                r_data[65] <= r_data[64];
                
                r_data[66] <= r_data[65];
                
                r_data[67] <= r_data[66];
                
                r_data[68] <= r_data[67];
                
                r_data[69] <= r_data[68];
                
                r_data[70] <= r_data[69];
                
                r_data[71] <= r_data[70];
                
                r_data[72] <= r_data[71];
                
                r_data[73] <= r_data[72];
                
                r_data[74] <= r_data[73];
                
                r_data[75] <= r_data[74];
                
                r_data[76] <= r_data[75];
                
                r_data[77] <= r_data[76];
                
                r_data[78] <= r_data[77];
                
                r_data[79] <= r_data[78];
                
                r_data[80] <= r_data[79];
                
                r_data[81] <= r_data[80];
                
                r_data[82] <= r_data[81];
                
                r_data[83] <= r_data[82];
                
                r_data[84] <= r_data[83];
                
                r_data[85] <= r_data[84];
                
                r_data[86] <= r_data[85];
                
                r_data[87] <= r_data[86];
                
                r_data[88] <= r_data[87];
                
                r_data[89] <= r_data[88];
                
                r_data[90] <= r_data[89];
                
                r_data[91] <= r_data[90];
                
                r_data[92] <= r_data[91];
                
                r_data[93] <= r_data[92];
                
                r_data[94] <= r_data[93];
                
                r_data[95] <= r_data[94];
                
                r_data[96] <= r_data[95];
                
                r_data[97] <= r_data[96];
                
                r_data[98] <= r_data[97];
                
                r_data[99] <= r_data[98];
                
                r_data[100] <= r_data[99];
                
                r_data[101] <= r_data[100];
                
                r_data[102] <= r_data[101];
                
                r_data[103] <= r_data[102];
                
                r_data[104] <= r_data[103];
                
                r_data[105] <= r_data[104];
                
                r_data[106] <= r_data[105];
                
                r_data[107] <= r_data[106];
                
                r_data[108] <= r_data[107];
                
                r_data[109] <= r_data[108];
                
                r_data[110] <= r_data[109];
                
                r_data[111] <= r_data[110];
                
                r_data[112] <= r_data[111];
                
                r_data[113] <= r_data[112];
                
                r_data[114] <= r_data[113];
                
                r_data[115] <= r_data[114];
                
                r_data[116] <= r_data[115];
                
                r_data[117] <= r_data[116];
                
                r_data[118] <= r_data[117];
                
                r_data[119] <= r_data[118];
                
                r_data[120] <= r_data[119];
                
                r_data[121] <= r_data[120];
                
                r_data[122] <= r_data[121];
                
                r_data[123] <= r_data[122];
                
                r_data[124] <= r_data[123];
                
                r_data[125] <= r_data[124];
                
                r_data[126] <= r_data[125];
                
                r_data[127] <= r_data[126];
                
                r_data[128] <= r_data[127];
                
                r_data[129] <= r_data[128];
                
                r_data[130] <= r_data[129];
                
                r_data[131] <= r_data[130];
                
                r_data[132] <= r_data[131];
                
                r_data[133] <= r_data[132];
                
                r_data[134] <= r_data[133];
                
                r_data[135] <= r_data[134];
                
                r_data[136] <= r_data[135];
                
                r_data[137] <= r_data[136];
                
                r_data[138] <= r_data[137];
                
                r_data[139] <= r_data[138];
                
                r_data[140] <= r_data[139];
                
                r_data[141] <= r_data[140];
                
                r_data[142] <= r_data[141];
                
                r_data[143] <= r_data[142];
                
                r_data[144] <= r_data[143];
                
                r_data[145] <= r_data[144];
                
                r_data[146] <= r_data[145];
                
                r_data[147] <= r_data[146];
                
                r_data[148] <= r_data[147];
                
                r_data[149] <= r_data[148];
                
                r_data[150] <= r_data[149];
                
                r_data[151] <= r_data[150];
                
                r_data[152] <= r_data[151];
                
                r_data[153] <= r_data[152];
                
                r_data[154] <= r_data[153];
                
                r_data[155] <= r_data[154];
                
                r_data[156] <= r_data[155];
                
                r_data[157] <= r_data[156];
                
                r_data[158] <= r_data[157];
                
                r_data[159] <= r_data[158];
                
                r_data[160] <= r_data[159];
                
                r_data[161] <= r_data[160];
                
                r_data[162] <= r_data[161];
                
                r_data[163] <= r_data[162];
                
                r_data[164] <= r_data[163];
                
                r_data[165] <= r_data[164];
                
                r_data[166] <= r_data[165];
                
                r_data[167] <= r_data[166];
                
                r_data[168] <= r_data[167];
                
                r_data[169] <= r_data[168];
                
                r_data[170] <= r_data[169];
                
                r_data[171] <= r_data[170];
                
                r_data[172] <= r_data[171];
                
                r_data[173] <= r_data[172];
                
                r_data[174] <= r_data[173];
                
                r_data[175] <= r_data[174];
                
                r_data[176] <= r_data[175];
                
                r_data[177] <= r_data[176];
                
                r_data[178] <= r_data[177];
                
                r_data[179] <= r_data[178];
                
                r_data[180] <= r_data[179];
                
                r_data[181] <= r_data[180];
                
                r_data[182] <= r_data[181];
                
                r_data[183] <= r_data[182];
                
                r_data[184] <= r_data[183];
                
                r_data[185] <= r_data[184];
                
                r_data[186] <= r_data[185];
                
                r_data[187] <= r_data[186];
                
                r_data[188] <= r_data[187];
                
                r_data[189] <= r_data[188];
                
                r_data[190] <= r_data[189];
                
                r_data[191] <= r_data[190];
                
                r_data[192] <= r_data[191];
                
                r_data[193] <= r_data[192];
                
                r_data[194] <= r_data[193];
                
                r_data[195] <= r_data[194];
                
                r_data[196] <= r_data[195];
                
                r_data[197] <= r_data[196];
                
                r_data[198] <= r_data[197];
                
                r_data[199] <= r_data[198];
                
                r_data[200] <= r_data[199];
                
                r_data[201] <= r_data[200];
                
                r_data[202] <= r_data[201];
                
                r_data[203] <= r_data[202];
                
                r_data[204] <= r_data[203];
                
                r_data[205] <= r_data[204];
                
                r_data[206] <= r_data[205];
                
                r_data[207] <= r_data[206];
                
                r_data[208] <= r_data[207];
                
                r_data[209] <= r_data[208];
                
                r_data[210] <= r_data[209];
                
                r_data[211] <= r_data[210];
                
                r_data[212] <= r_data[211];
                
                r_data[213] <= r_data[212];
                
                r_data[214] <= r_data[213];
                
                r_data[215] <= r_data[214];
                
                r_data[216] <= r_data[215];
                
                r_data[217] <= r_data[216];
                
                r_data[218] <= r_data[217];
                
                r_data[219] <= r_data[218];
                
                r_data[220] <= r_data[219];
                
                r_data[221] <= r_data[220];
                
                r_data[222] <= r_data[221];
                
                r_data[223] <= r_data[222];
                
                r_data[224] <= r_data[223];
                
                r_data[225] <= r_data[224];
                
                r_data[226] <= r_data[225];
                
                r_data[227] <= r_data[226];
                
                r_data[228] <= r_data[227];
                
                r_data[229] <= r_data[228];
                
                r_data[230] <= r_data[229];
                
                r_data[231] <= r_data[230];
                
                r_data[232] <= r_data[231];
                
                r_data[233] <= r_data[232];
                
                r_data[234] <= r_data[233];
                
                r_data[235] <= r_data[234];
                
                r_data[236] <= r_data[235];
                
                r_data[237] <= r_data[236];
                
                r_data[238] <= r_data[237];
                
                r_data[239] <= r_data[238];
                
                r_data[240] <= r_data[239];
                
                r_data[241] <= r_data[240];
                
                r_data[242] <= r_data[241];
                
                r_data[243] <= r_data[242];
                
                r_data[244] <= r_data[243];
                
                r_data[245] <= r_data[244];
                
                r_data[246] <= r_data[245];
                
                r_data[247] <= r_data[246];
                
                r_data[248] <= r_data[247];
                
                r_data[249] <= r_data[248];
                
                r_data[250] <= r_data[249];
                
                r_data[251] <= r_data[250];
                
                r_data[252] <= r_data[251];
                
                r_data[253] <= r_data[252];
                
                r_data[254] <= r_data[253];
                
                r_data[255] <= r_data[254];
                
                r_data[256] <= r_data[255];
                
                r_data[257] <= r_data[256];
                
                r_data[258] <= r_data[257];
                
                r_data[259] <= r_data[258];
                
                r_data[260] <= r_data[259];
                
                r_data[261] <= r_data[260];
                
                r_data[262] <= r_data[261];
                
                r_data[263] <= r_data[262];
                
                r_data[264] <= r_data[263];
                
                r_data[265] <= r_data[264];
                
                r_data[266] <= r_data[265];
                
                r_data[267] <= r_data[266];
                
                r_data[268] <= r_data[267];
                
                r_data[269] <= r_data[268];
                
                r_data[270] <= r_data[269];
                
                r_data[271] <= r_data[270];
                
                r_data[272] <= r_data[271];
                
                r_data[273] <= r_data[272];
                
                r_data[274] <= r_data[273];
                
                r_data[275] <= r_data[274];
                
                r_data[276] <= r_data[275];
                
                r_data[277] <= r_data[276];
                
                r_data[278] <= r_data[277];
                
                r_data[279] <= r_data[278];
                
                r_data[280] <= r_data[279];
                
                r_data[281] <= r_data[280];
                
                r_data[282] <= r_data[281];
                
                r_data[283] <= r_data[282];
                
                r_data[284] <= r_data[283];
                
                r_data[285] <= r_data[284];
                
                r_data[286] <= r_data[285];
                
                r_data[287] <= r_data[286];
                
                r_data[288] <= r_data[287];
                
                r_data[289] <= r_data[288];
                
                r_data[290] <= r_data[289];
                
                r_data[291] <= r_data[290];
                
                r_data[292] <= r_data[291];
                
                r_data[293] <= r_data[292];
                
                r_data[294] <= r_data[293];
                
                r_data[295] <= r_data[294];
                
                r_data[296] <= r_data[295];
                
                r_data[297] <= r_data[296];
                
                r_data[298] <= r_data[297];
                
                r_data[299] <= r_data[298];
                
                r_data[300] <= r_data[299];
                
                r_data[301] <= r_data[300];
                
                r_data[302] <= r_data[301];
                
                r_data[303] <= r_data[302];
                
                r_data[304] <= r_data[303];
                
                r_data[305] <= r_data[304];
                
                r_data[306] <= r_data[305];
                
                r_data[307] <= r_data[306];
                
                r_data[308] <= r_data[307];
                
                r_data[309] <= r_data[308];
                
                r_data[310] <= r_data[309];
                
                r_data[311] <= r_data[310];
                
                r_data[312] <= r_data[311];
                
                r_data[313] <= r_data[312];
                
                r_data[314] <= r_data[313];
                
                r_data[315] <= r_data[314];
                
                r_data[316] <= r_data[315];
                
                r_data[317] <= r_data[316];
                
                r_data[318] <= r_data[317];
                
                r_data[319] <= r_data[318];
                
                r_data[320] <= r_data[319];
                
                r_data[321] <= r_data[320];
                
                r_data[322] <= r_data[321];
                
                r_data[323] <= r_data[322];
                
                r_data[324] <= r_data[323];
                
                r_data[325] <= r_data[324];
                
                r_data[326] <= r_data[325];
                
                r_data[327] <= r_data[326];
                
                r_data[328] <= r_data[327];
                
                r_data[329] <= r_data[328];
                
                r_data[330] <= r_data[329];
                
                r_data[331] <= r_data[330];
                
                r_data[332] <= r_data[331];
                
                r_data[333] <= r_data[332];
                
                r_data[334] <= r_data[333];
                
                r_data[335] <= r_data[334];
                
                r_data[336] <= r_data[335];
                
                r_data[337] <= r_data[336];
                
                r_data[338] <= r_data[337];
                
                r_data[339] <= r_data[338];
                
                r_data[340] <= r_data[339];
                
                r_data[341] <= r_data[340];
                
                r_data[342] <= r_data[341];
                
                r_data[343] <= r_data[342];
                
                r_data[344] <= r_data[343];
                
                r_data[345] <= r_data[344];
                
                r_data[346] <= r_data[345];
                
                r_data[347] <= r_data[346];
                
                r_data[348] <= r_data[347];
                
                r_data[349] <= r_data[348];
                
                r_data[350] <= r_data[349];
                
                r_data[351] <= r_data[350];
                
                r_data[352] <= r_data[351];
                
                r_data[353] <= r_data[352];
                
                r_data[354] <= r_data[353];
                
                r_data[355] <= r_data[354];
                
                r_data[356] <= r_data[355];
                
                r_data[357] <= r_data[356];
                
                r_data[358] <= r_data[357];
                
                r_data[359] <= r_data[358];
                
                r_data[360] <= r_data[359];
                
                r_data[361] <= r_data[360];
                
                r_data[362] <= r_data[361];
                
                r_data[363] <= r_data[362];
                
                r_data[364] <= r_data[363];
                
                r_data[365] <= r_data[364];
                
                r_data[366] <= r_data[365];
                
                r_data[367] <= r_data[366];
                
                r_data[368] <= r_data[367];
                
                r_data[369] <= r_data[368];
                
                r_data[370] <= r_data[369];
                
                r_data[371] <= r_data[370];
                
                r_data[372] <= r_data[371];
                
                r_data[373] <= r_data[372];
                
                r_data[374] <= r_data[373];
                
                r_data[375] <= r_data[374];
                
                r_data[376] <= r_data[375];
                
                r_data[377] <= r_data[376];
                
                r_data[378] <= r_data[377];
                
                r_data[379] <= r_data[378];
                
                r_data[380] <= r_data[379];
                
                r_data[381] <= r_data[380];
                
                r_data[382] <= r_data[381];
                
                r_data[383] <= r_data[382];
                
                r_data[384] <= r_data[383];
                
                r_data[385] <= r_data[384];
                
                r_data[386] <= r_data[385];
                
                r_data[387] <= r_data[386];
                
                r_data[388] <= r_data[387];
                
                r_data[389] <= r_data[388];
                
                r_data[390] <= r_data[389];
                
                r_data[391] <= r_data[390];
                
                r_data[392] <= r_data[391];
                
                r_data[393] <= r_data[392];
                
                r_data[394] <= r_data[393];
                
                r_data[395] <= r_data[394];
                
                r_data[396] <= r_data[395];
                
                r_data[397] <= r_data[396];
                
                r_data[398] <= r_data[397];
                
                r_data[399] <= r_data[398];
                
                r_data[400] <= r_data[399];
                
                r_data[401] <= r_data[400];
                
                r_data[402] <= r_data[401];
                
                r_data[403] <= r_data[402];
                
                r_data[404] <= r_data[403];
                
                r_data[405] <= r_data[404];
                
                r_data[406] <= r_data[405];
                
                r_data[407] <= r_data[406];
                
                r_data[408] <= r_data[407];
                
                r_data[409] <= r_data[408];
                
                r_data[410] <= r_data[409];
                
                r_data[411] <= r_data[410];
                
                r_data[412] <= r_data[411];
                
                r_data[413] <= r_data[412];
                
                r_data[414] <= r_data[413];
                
                r_data[415] <= r_data[414];
                
                r_data[416] <= r_data[415];
                
                r_data[417] <= r_data[416];
                
                r_data[418] <= r_data[417];
                
                r_data[419] <= r_data[418];
                
                r_data[420] <= r_data[419];
                
                r_data[421] <= r_data[420];
                
                r_data[422] <= r_data[421];
                
                r_data[423] <= r_data[422];
                
                r_data[424] <= r_data[423];
                
                r_data[425] <= r_data[424];
                
                r_data[426] <= r_data[425];
                
                r_data[427] <= r_data[426];
                
                r_data[428] <= r_data[427];
                
                r_data[429] <= r_data[428];
                
                r_data[430] <= r_data[429];
                
                r_data[431] <= r_data[430];
                
                r_data[432] <= r_data[431];
                
                r_data[433] <= r_data[432];
                
                r_data[434] <= r_data[433];
                
                r_data[435] <= r_data[434];
                
                r_data[436] <= r_data[435];
                
                r_data[437] <= r_data[436];
                
                r_data[438] <= r_data[437];
                
                r_data[439] <= r_data[438];
                
                r_data[440] <= r_data[439];
                
                r_data[441] <= r_data[440];
                
                r_data[442] <= r_data[441];
                
                r_data[443] <= r_data[442];
                
                r_data[444] <= r_data[443];
                
                r_data[445] <= r_data[444];
                
                r_data[446] <= r_data[445];
                
                r_data[447] <= r_data[446];
                
                r_data[448] <= r_data[447];
                
                r_data[449] <= r_data[448];
                
                r_data[450] <= r_data[449];
                
                r_data[451] <= r_data[450];
                
                r_data[452] <= r_data[451];
                
                r_data[453] <= r_data[452];
                
                r_data[454] <= r_data[453];
                
                r_data[455] <= r_data[454];
                
                r_data[456] <= r_data[455];
                
                r_data[457] <= r_data[456];
                
                r_data[458] <= r_data[457];
                
                r_data[459] <= r_data[458];
                
                r_data[460] <= r_data[459];
                
                r_data[461] <= r_data[460];
                
                r_data[462] <= r_data[461];
                
                r_data[463] <= r_data[462];
                
                r_data[464] <= r_data[463];
                
                r_data[465] <= r_data[464];
                
                r_data[466] <= r_data[465];
                
                r_data[467] <= r_data[466];
                
                r_data[468] <= r_data[467];
                
                r_data[469] <= r_data[468];
                
                r_data[470] <= r_data[469];
                
                r_data[471] <= r_data[470];
                
                r_data[472] <= r_data[471];
                
                r_data[473] <= r_data[472];
                
                r_data[474] <= r_data[473];
                
                r_data[475] <= r_data[474];
                
                r_data[476] <= r_data[475];
                
                r_data[477] <= r_data[476];
                
                r_data[478] <= r_data[477];
                
                r_data[479] <= r_data[478];
                
                r_data[480] <= r_data[479];
                
                r_data[481] <= r_data[480];
                
                r_data[482] <= r_data[481];
                
                r_data[483] <= r_data[482];
                
                r_data[484] <= r_data[483];
                
                r_data[485] <= r_data[484];
                
                r_data[486] <= r_data[485];
                
                r_data[487] <= r_data[486];
                
                r_data[488] <= r_data[487];
                
                r_data[489] <= r_data[488];
                
                r_data[490] <= r_data[489];
                
                r_data[491] <= r_data[490];
                
                r_data[492] <= r_data[491];
                
                r_data[493] <= r_data[492];
                
                r_data[494] <= r_data[493];
                
                r_data[495] <= r_data[494];
                
                r_data[496] <= r_data[495];
                
                r_data[497] <= r_data[496];
                
                r_data[498] <= r_data[497];
                
                r_data[499] <= r_data[498];
                
                r_data[500] <= r_data[499];
                
                r_data[501] <= r_data[500];
                
                r_data[502] <= r_data[501];
                
                r_data[503] <= r_data[502];
                
                r_data[504] <= r_data[503];
                
                r_data[505] <= r_data[504];
                
                r_data[506] <= r_data[505];
                
                r_data[507] <= r_data[506];
                
                r_data[508] <= r_data[507];
                
                r_data[509] <= r_data[508];
                
                r_data[510] <= r_data[509];
                
                r_data[511] <= r_data[510];
                
                r_data[512] <= r_data[511];
                
                r_data[513] <= r_data[512];
                
                r_data[514] <= r_data[513];
                
                r_data[515] <= r_data[514];
                
                r_data[516] <= r_data[515];
                
                r_data[517] <= r_data[516];
                
                r_data[518] <= r_data[517];
                
                r_data[519] <= r_data[518];
                
                r_data[520] <= r_data[519];
                
                r_data[521] <= r_data[520];
                
                r_data[522] <= r_data[521];
                
                r_data[523] <= r_data[522];
                
                r_data[524] <= r_data[523];
                
                r_data[525] <= r_data[524];
                
                r_data[526] <= r_data[525];
                
                r_data[527] <= r_data[526];
                
                r_data[528] <= r_data[527];
                
                r_data[529] <= r_data[528];
                
                r_data[530] <= r_data[529];
                
                r_data[531] <= r_data[530];
                
                r_data[532] <= r_data[531];
                
                r_data[533] <= r_data[532];
                
                r_data[534] <= r_data[533];
                
                r_data[535] <= r_data[534];
                
                r_data[536] <= r_data[535];
                
                r_data[537] <= r_data[536];
                
                r_data[538] <= r_data[537];
                
                r_data[539] <= r_data[538];
                
                r_data[540] <= r_data[539];
                
                r_data[541] <= r_data[540];
                
                r_data[542] <= r_data[541];
                
                r_data[543] <= r_data[542];
                
                r_data[544] <= r_data[543];
                
                r_data[545] <= r_data[544];
                
                r_data[546] <= r_data[545];
                
                r_data[547] <= r_data[546];
                
                r_data[548] <= r_data[547];
                
                r_data[549] <= r_data[548];
                
                r_data[550] <= r_data[549];
                
                r_data[551] <= r_data[550];
                
                r_data[552] <= r_data[551];
                
                r_data[553] <= r_data[552];
                
                r_data[554] <= r_data[553];
                
                r_data[555] <= r_data[554];
                
                r_data[556] <= r_data[555];
                
                r_data[557] <= r_data[556];
                
                r_data[558] <= r_data[557];
                
                r_data[559] <= r_data[558];
                
                r_data[560] <= r_data[559];
                
                r_data[561] <= r_data[560];
                
                r_data[562] <= r_data[561];
                
                r_data[563] <= r_data[562];
                
                r_data[564] <= r_data[563];
                
                r_data[565] <= r_data[564];
                
                r_data[566] <= r_data[565];
                
                r_data[567] <= r_data[566];
                
                r_data[568] <= r_data[567];
                
                r_data[569] <= r_data[568];
                
                r_data[570] <= r_data[569];
                
                r_data[571] <= r_data[570];
                
                r_data[572] <= r_data[571];
                
                r_data[573] <= r_data[572];
                
                r_data[574] <= r_data[573];
                
                r_data[575] <= r_data[574];
                
                r_data[576] <= r_data[575];
                
                r_data[577] <= r_data[576];
                
                r_data[578] <= r_data[577];
                
                r_data[579] <= r_data[578];
                
                r_data[580] <= r_data[579];
                
                r_data[581] <= r_data[580];
                
                r_data[582] <= r_data[581];
                
                r_data[583] <= r_data[582];
                
                r_data[584] <= r_data[583];
                
                r_data[585] <= r_data[584];
                
                r_data[586] <= r_data[585];
                
                r_data[587] <= r_data[586];
                
                r_data[588] <= r_data[587];
                
                r_data[589] <= r_data[588];
                
                r_data[590] <= r_data[589];
                
                r_data[591] <= r_data[590];
                
                r_data[592] <= r_data[591];
                
                r_data[593] <= r_data[592];
                
                r_data[594] <= r_data[593];
                
                r_data[595] <= r_data[594];
                
                r_data[596] <= r_data[595];
                
                r_data[597] <= r_data[596];
                
                r_data[598] <= r_data[597];
                
                r_data[599] <= r_data[598];
                
                r_data[600] <= r_data[599];
                
                r_data[601] <= r_data[600];
                
                r_data[602] <= r_data[601];
                
                r_data[603] <= r_data[602];
                
                r_data[604] <= r_data[603];
                
                r_data[605] <= r_data[604];
                
                r_data[606] <= r_data[605];
                
                r_data[607] <= r_data[606];
                
                r_data[608] <= r_data[607];
                
                r_data[609] <= r_data[608];
                
                r_data[610] <= r_data[609];
                
                r_data[611] <= r_data[610];
                
                r_data[612] <= r_data[611];
                
                r_data[613] <= r_data[612];
                
                r_data[614] <= r_data[613];
                
                r_data[615] <= r_data[614];
                
                r_data[616] <= r_data[615];
                
                r_data[617] <= r_data[616];
                
                r_data[618] <= r_data[617];
                
                r_data[619] <= r_data[618];
                
                r_data[620] <= r_data[619];
                
                r_data[621] <= r_data[620];
                
                r_data[622] <= r_data[621];
                
                r_data[623] <= r_data[622];
                
                r_data[624] <= r_data[623];
                
                r_data[625] <= r_data[624];
                
                r_data[626] <= r_data[625];
                
                r_data[627] <= r_data[626];
                
                r_data[628] <= r_data[627];
                
                r_data[629] <= r_data[628];
                
                r_data[630] <= r_data[629];
                
                r_data[631] <= r_data[630];
                
                r_data[632] <= r_data[631];
                
                r_data[633] <= r_data[632];
                
                r_data[634] <= r_data[633];
                
                r_data[635] <= r_data[634];
                
                r_data[636] <= r_data[635];
                
                r_data[637] <= r_data[636];
                
                r_data[638] <= r_data[637];
                
                r_data[639] <= r_data[638];
                
                r_data[640] <= r_data[639];
                
                r_data[641] <= r_data[640];
                
                r_data[642] <= r_data[641];
                
                r_data[643] <= r_data[642];
                
                r_data[644] <= r_data[643];
                
                r_data[645] <= r_data[644];
                
                r_data[646] <= r_data[645];
                
                r_data[647] <= r_data[646];
                
                r_data[648] <= r_data[647];
                
                r_data[649] <= r_data[648];
                
                r_data[650] <= r_data[649];
                
                r_data[651] <= r_data[650];
                
                r_data[652] <= r_data[651];
                
                r_data[653] <= r_data[652];
                
                r_data[654] <= r_data[653];
                
                r_data[655] <= r_data[654];
                
                r_data[656] <= r_data[655];
                
                r_data[657] <= r_data[656];
                
                r_data[658] <= r_data[657];
                
                r_data[659] <= r_data[658];
                
                r_data[660] <= r_data[659];
                
                r_data[661] <= r_data[660];
                
                r_data[662] <= r_data[661];
                
                r_data[663] <= r_data[662];
                
                r_data[664] <= r_data[663];
                
                r_data[665] <= r_data[664];
                
                r_data[666] <= r_data[665];
                
                r_data[667] <= r_data[666];
                
                r_data[668] <= r_data[667];
                
                r_data[669] <= r_data[668];
                
                r_data[670] <= r_data[669];
                
                r_data[671] <= r_data[670];
                
                r_data[672] <= r_data[671];
                
                r_data[673] <= r_data[672];
                
                r_data[674] <= r_data[673];
                
                r_data[675] <= r_data[674];
                
                r_data[676] <= r_data[675];
                
                r_data[677] <= r_data[676];
                
                r_data[678] <= r_data[677];
                
                r_data[679] <= r_data[678];
                
                r_data[680] <= r_data[679];
                
                r_data[681] <= r_data[680];
                
                r_data[682] <= r_data[681];
                
                r_data[683] <= r_data[682];
                
                r_data[684] <= r_data[683];
                
                r_data[685] <= r_data[684];
                
                r_data[686] <= r_data[685];
                
                r_data[687] <= r_data[686];
                
                r_data[688] <= r_data[687];
                
                r_data[689] <= r_data[688];
                
                r_data[690] <= r_data[689];
                
                r_data[691] <= r_data[690];
                
                r_data[692] <= r_data[691];
                
                r_data[693] <= r_data[692];
                
                r_data[694] <= r_data[693];
                
                r_data[695] <= r_data[694];
                
                r_data[696] <= r_data[695];
                
                r_data[697] <= r_data[696];
                
                r_data[698] <= r_data[697];
                
                r_data[699] <= r_data[698];
                
                r_data[700] <= r_data[699];
                
                r_data[701] <= r_data[700];
                
                r_data[702] <= r_data[701];
                
                r_data[703] <= r_data[702];
                
                r_data[704] <= r_data[703];
                
                r_data[705] <= r_data[704];
                
                r_data[706] <= r_data[705];
                
                r_data[707] <= r_data[706];
                
                r_data[708] <= r_data[707];
                
                r_data[709] <= r_data[708];
                
                r_data[710] <= r_data[709];
                
                r_data[711] <= r_data[710];
                
                r_data[712] <= r_data[711];
                
                r_data[713] <= r_data[712];
                
                r_data[714] <= r_data[713];
                
                r_data[715] <= r_data[714];
                
                r_data[716] <= r_data[715];
                
                r_data[717] <= r_data[716];
                
                r_data[718] <= r_data[717];
                
                r_data[719] <= r_data[718];
                
                r_data[720] <= r_data[719];
                
                r_data[721] <= r_data[720];
                
                r_data[722] <= r_data[721];
                
                r_data[723] <= r_data[722];
                
                r_data[724] <= r_data[723];
                
                r_data[725] <= r_data[724];
                
                r_data[726] <= r_data[725];
                
                r_data[727] <= r_data[726];
                
                r_data[728] <= r_data[727];
                
                r_data[729] <= r_data[728];
                
                r_data[730] <= r_data[729];
                
                r_data[731] <= r_data[730];
                
                r_data[732] <= r_data[731];
                
                r_data[733] <= r_data[732];
                
                r_data[734] <= r_data[733];
                
                r_data[735] <= r_data[734];
                
                r_data[736] <= r_data[735];
                
                r_data[737] <= r_data[736];
                
                r_data[738] <= r_data[737];
                
                r_data[739] <= r_data[738];
                
                r_data[740] <= r_data[739];
                
                r_data[741] <= r_data[740];
                
                r_data[742] <= r_data[741];
                
                r_data[743] <= r_data[742];
                
                r_data[744] <= r_data[743];
                
                r_data[745] <= r_data[744];
                
                r_data[746] <= r_data[745];
                
                r_data[747] <= r_data[746];
                
                r_data[748] <= r_data[747];
                
                r_data[749] <= r_data[748];
                
                r_data[750] <= r_data[749];
                
                r_data[751] <= r_data[750];
                
                r_data[752] <= r_data[751];
                
                r_data[753] <= r_data[752];
                
                r_data[754] <= r_data[753];
                
                r_data[755] <= r_data[754];
                
                r_data[756] <= r_data[755];
                
                r_data[757] <= r_data[756];
                
                r_data[758] <= r_data[757];
                
                r_data[759] <= r_data[758];
                
                r_data[760] <= r_data[759];
                
                r_data[761] <= r_data[760];
                
                r_data[762] <= r_data[761];
                
                r_data[763] <= r_data[762];
                
                r_data[764] <= r_data[763];
                
                r_data[765] <= r_data[764];
                
                r_data[766] <= r_data[765];
                
                r_data[767] <= r_data[766];
                
                r_data[768] <= r_data[767];
                
                r_data[769] <= r_data[768];
                
                r_data[770] <= r_data[769];
                
                r_data[771] <= r_data[770];
                
                r_data[772] <= r_data[771];
                
                r_data[773] <= r_data[772];
                
                r_data[774] <= r_data[773];
                
                r_data[775] <= r_data[774];
                
                r_data[776] <= r_data[775];
                
                r_data[777] <= r_data[776];
                
                r_data[778] <= r_data[777];
                
                r_data[779] <= r_data[778];
                
                r_data[780] <= r_data[779];
                
                r_data[781] <= r_data[780];
                
                r_data[782] <= r_data[781];
                
                r_data[783] <= r_data[782];
                
                r_data[784] <= r_data[783];
                
                r_data[785] <= r_data[784];
                
                r_data[786] <= r_data[785];
                
                r_data[787] <= r_data[786];
                
                r_data[788] <= r_data[787];
                
                r_data[789] <= r_data[788];
                
                r_data[790] <= r_data[789];
                
                r_data[791] <= r_data[790];
                
                r_data[792] <= r_data[791];
                
                r_data[793] <= r_data[792];
                
                r_data[794] <= r_data[793];
                
                r_data[795] <= r_data[794];
                
                r_data[796] <= r_data[795];
                
                r_data[797] <= r_data[796];
                
                r_data[798] <= r_data[797];
                
                r_data[799] <= r_data[798];
                
                r_data[800] <= r_data[799];
                
                r_data[801] <= r_data[800];
                
                r_data[802] <= r_data[801];
                
                r_data[803] <= r_data[802];
                
                r_data[804] <= r_data[803];
                
                r_data[805] <= r_data[804];
                
                r_data[806] <= r_data[805];
                
                r_data[807] <= r_data[806];
                
                r_data[808] <= r_data[807];
                
                r_data[809] <= r_data[808];
                
                r_data[810] <= r_data[809];
                
                r_data[811] <= r_data[810];
                
                r_data[812] <= r_data[811];
                
                r_data[813] <= r_data[812];
                
                r_data[814] <= r_data[813];
                
                r_data[815] <= r_data[814];
                
                r_data[816] <= r_data[815];
                
                r_data[817] <= r_data[816];
                
                r_data[818] <= r_data[817];
                
                r_data[819] <= r_data[818];
                
                r_data[820] <= r_data[819];
                
                r_data[821] <= r_data[820];
                
                r_data[822] <= r_data[821];
                
                r_data[823] <= r_data[822];
                
                r_data[824] <= r_data[823];
                
                r_data[825] <= r_data[824];
                
                r_data[826] <= r_data[825];
                
                r_data[827] <= r_data[826];
                
                r_data[828] <= r_data[827];
                
                r_data[829] <= r_data[828];
                
                r_data[830] <= r_data[829];
                
                r_data[831] <= r_data[830];
                
                r_data[832] <= r_data[831];
                
                r_data[833] <= r_data[832];
                
                r_data[834] <= r_data[833];
                
                r_data[835] <= r_data[834];
                
                r_data[836] <= r_data[835];
                
                r_data[837] <= r_data[836];
                
                r_data[838] <= r_data[837];
                
                r_data[839] <= r_data[838];
                
                r_data[840] <= r_data[839];
                
                r_data[841] <= r_data[840];
                
                r_data[842] <= r_data[841];
                
                r_data[843] <= r_data[842];
                
                r_data[844] <= r_data[843];
                
                r_data[845] <= r_data[844];
                
                r_data[846] <= r_data[845];
                
                r_data[847] <= r_data[846];
                
                r_data[848] <= r_data[847];
                
                r_data[849] <= r_data[848];
                
                r_data[850] <= r_data[849];
                
                r_data[851] <= r_data[850];
                
                r_data[852] <= r_data[851];
                
                r_data[853] <= r_data[852];
                
                r_data[854] <= r_data[853];
                
                r_data[855] <= r_data[854];
                
                r_data[856] <= r_data[855];
                
                r_data[857] <= r_data[856];
                
                r_data[858] <= r_data[857];
                
                r_data[859] <= r_data[858];
                
                r_data[860] <= r_data[859];
                
                r_data[861] <= r_data[860];
                
                r_data[862] <= r_data[861];
                
                r_data[863] <= r_data[862];
                
                r_data[864] <= r_data[863];
                
                r_data[865] <= r_data[864];
                
                r_data[866] <= r_data[865];
                
                r_data[867] <= r_data[866];
                
                r_data[868] <= r_data[867];
                
                r_data[869] <= r_data[868];
                
                r_data[870] <= r_data[869];
                
                r_data[871] <= r_data[870];
                
                r_data[872] <= r_data[871];
                
                r_data[873] <= r_data[872];
                
                r_data[874] <= r_data[873];
                
                r_data[875] <= r_data[874];
                
                r_data[876] <= r_data[875];
                
                r_data[877] <= r_data[876];
                
                r_data[878] <= r_data[877];
                
                r_data[879] <= r_data[878];
                
                r_data[880] <= r_data[879];
                
                r_data[881] <= r_data[880];
                
                r_data[882] <= r_data[881];
                
                r_data[883] <= r_data[882];
                
                r_data[884] <= r_data[883];
                
                r_data[885] <= r_data[884];
                
                r_data[886] <= r_data[885];
                
                r_data[887] <= r_data[886];
                
                r_data[888] <= r_data[887];
                
                r_data[889] <= r_data[888];
                
                r_data[890] <= r_data[889];
                
                r_data[891] <= r_data[890];
                
                r_data[892] <= r_data[891];
                
                r_data[893] <= r_data[892];
                
                r_data[894] <= r_data[893];
                
                r_data[895] <= r_data[894];
                
                r_data[896] <= r_data[895];
                
                r_data[897] <= r_data[896];
                
                r_data[898] <= r_data[897];
                
                r_data[899] <= r_data[898];
                
                r_data[900] <= r_data[899];
                
                r_data[901] <= r_data[900];
                
                r_data[902] <= r_data[901];
                
                r_data[903] <= r_data[902];
                
                r_data[904] <= r_data[903];
                
                r_data[905] <= r_data[904];
                
                r_data[906] <= r_data[905];
                
                r_data[907] <= r_data[906];
                
                r_data[908] <= r_data[907];
                
                r_data[909] <= r_data[908];
                
                r_data[910] <= r_data[909];
                
                r_data[911] <= r_data[910];
                
                r_data[912] <= r_data[911];
                
                r_data[913] <= r_data[912];
                
                r_data[914] <= r_data[913];
                
                r_data[915] <= r_data[914];
                
                r_data[916] <= r_data[915];
                
                r_data[917] <= r_data[916];
                
                r_data[918] <= r_data[917];
                
                r_data[919] <= r_data[918];
                
                r_data[920] <= r_data[919];
                
                r_data[921] <= r_data[920];
                
                r_data[922] <= r_data[921];
                
                r_data[923] <= r_data[922];
                
                r_data[924] <= r_data[923];
                
                r_data[925] <= r_data[924];
                
                r_data[926] <= r_data[925];
                
                r_data[927] <= r_data[926];
                
                r_data[928] <= r_data[927];
                
                r_data[929] <= r_data[928];
                
                r_data[930] <= r_data[929];
                
                r_data[931] <= r_data[930];
                
                r_data[932] <= r_data[931];
                
                r_data[933] <= r_data[932];
                
                r_data[934] <= r_data[933];
                
                r_data[935] <= r_data[934];
                
                r_data[936] <= r_data[935];
                
                r_data[937] <= r_data[936];
                
                r_data[938] <= r_data[937];
                
                r_data[939] <= r_data[938];
                
                r_data[940] <= r_data[939];
                
                r_data[941] <= r_data[940];
                
                r_data[942] <= r_data[941];
                
                r_data[943] <= r_data[942];
                
                r_data[944] <= r_data[943];
                
                r_data[945] <= r_data[944];
                
                r_data[946] <= r_data[945];
                
                r_data[947] <= r_data[946];
                
                r_data[948] <= r_data[947];
                
                r_data[949] <= r_data[948];
                
                r_data[950] <= r_data[949];
                
                r_data[951] <= r_data[950];
                
                r_data[952] <= r_data[951];
                
                r_data[953] <= r_data[952];
                
                r_data[954] <= r_data[953];
                
                r_data[955] <= r_data[954];
                
                r_data[956] <= r_data[955];
                
                r_data[957] <= r_data[956];
                
                r_data[958] <= r_data[957];
                
                r_data[959] <= r_data[958];
                
                r_data[960] <= r_data[959];
                
                r_data[961] <= r_data[960];
                
                r_data[962] <= r_data[961];
                
                r_data[963] <= r_data[962];
                
                r_data[964] <= r_data[963];
                
                r_data[965] <= r_data[964];
                
                r_data[966] <= r_data[965];
                
                r_data[967] <= r_data[966];
                
                r_data[968] <= r_data[967];
                
                r_data[969] <= r_data[968];
                
                r_data[970] <= r_data[969];
                
                r_data[971] <= r_data[970];
                
                r_data[972] <= r_data[971];
                
                r_data[973] <= r_data[972];
                
                r_data[974] <= r_data[973];
                
                r_data[975] <= r_data[974];
                
                r_data[976] <= r_data[975];
                
                r_data[977] <= r_data[976];
                
                r_data[978] <= r_data[977];
                
                r_data[979] <= r_data[978];
                
                r_data[980] <= r_data[979];
                
                r_data[981] <= r_data[980];
                
                r_data[982] <= r_data[981];
                
                r_data[983] <= r_data[982];
                
                r_data[984] <= r_data[983];
                
                r_data[985] <= r_data[984];
                
                r_data[986] <= r_data[985];
                
                r_data[987] <= r_data[986];
                
                r_data[988] <= r_data[987];
                
                r_data[989] <= r_data[988];
                
                r_data[990] <= r_data[989];
                
                r_data[991] <= r_data[990];
                
                r_data[992] <= r_data[991];
                
                r_data[993] <= r_data[992];
                
                r_data[994] <= r_data[993];
                
                r_data[995] <= r_data[994];
                
                r_data[996] <= r_data[995];
                
                r_data[997] <= r_data[996];
                
                r_data[998] <= r_data[997];
                
                r_data[999] <= r_data[998];
                
                r_data[1000] <= r_data[999];
                
                r_data[1001] <= r_data[1000];
                
                r_data[1002] <= r_data[1001];
                
                r_data[1003] <= r_data[1002];
                
                r_data[1004] <= r_data[1003];
                
                r_data[1005] <= r_data[1004];
                
                r_data[1006] <= r_data[1005];
                
                r_data[1007] <= r_data[1006];
                
                r_data[1008] <= r_data[1007];
                
                r_data[1009] <= r_data[1008];
                
                r_data[1010] <= r_data[1009];
                
                r_data[1011] <= r_data[1010];
                
                r_data[1012] <= r_data[1011];
                
                r_data[1013] <= r_data[1012];
                
                r_data[1014] <= r_data[1013];
                
                r_data[1015] <= r_data[1014];
                
                r_data[1016] <= r_data[1015];
                
                r_data[1017] <= r_data[1016];
                
                r_data[1018] <= r_data[1017];
                
                r_data[1019] <= r_data[1018];
                
                r_data[1020] <= r_data[1019];
                
                r_data[1021] <= r_data[1020];
                
                r_data[1022] <= r_data[1021];
                
                r_data[1023] <= r_data[1022];
                
                r_data[1024] <= r_data[1023];
                
                r_data[1025] <= r_data[1024];
                
                r_data[1026] <= r_data[1025];
                
                r_data[1027] <= r_data[1026];
                
                r_data[1028] <= r_data[1027];
                
                r_data[1029] <= r_data[1028];
                
                r_data[1030] <= r_data[1029];
                
                r_data[1031] <= r_data[1030];
                
                r_data[1032] <= r_data[1031];
                
                r_data[1033] <= r_data[1032];
                
                r_data[1034] <= r_data[1033];
                
                r_data[1035] <= r_data[1034];
                
                r_data[1036] <= r_data[1035];
                
                r_data[1037] <= r_data[1036];
                
                r_data[1038] <= r_data[1037];
                
                r_data[1039] <= r_data[1038];
                
                r_data[1040] <= r_data[1039];
                
                r_data[1041] <= r_data[1040];
                
                r_data[1042] <= r_data[1041];
                
                r_data[1043] <= r_data[1042];
                
                r_data[1044] <= r_data[1043];
                
                r_data[1045] <= r_data[1044];
                
                r_data[1046] <= r_data[1045];
                
                r_data[1047] <= r_data[1046];
                
                r_data[1048] <= r_data[1047];
                
                r_data[1049] <= r_data[1048];
                
                r_data[1050] <= r_data[1049];
                
                r_data[1051] <= r_data[1050];
                
                r_data[1052] <= r_data[1051];
                
                r_data[1053] <= r_data[1052];
                
                r_data[1054] <= r_data[1053];
                
                r_data[1055] <= r_data[1054];
                
                r_data[1056] <= r_data[1055];
                
                r_data[1057] <= r_data[1056];
                
                r_data[1058] <= r_data[1057];
                
                r_data[1059] <= r_data[1058];
                
                r_data[1060] <= r_data[1059];
                
                r_data[1061] <= r_data[1060];
                
                r_data[1062] <= r_data[1061];
                
                r_data[1063] <= r_data[1062];
                
                r_data[1064] <= r_data[1063];
                
                r_data[1065] <= r_data[1064];
                
                r_data[1066] <= r_data[1065];
                
                r_data[1067] <= r_data[1066];
                
                r_data[1068] <= r_data[1067];
                
                r_data[1069] <= r_data[1068];
                
                r_data[1070] <= r_data[1069];
                
                r_data[1071] <= r_data[1070];
                
                r_data[1072] <= r_data[1071];
                
                r_data[1073] <= r_data[1072];
                
                r_data[1074] <= r_data[1073];
                
                r_data[1075] <= r_data[1074];
                
                r_data[1076] <= r_data[1075];
                
                r_data[1077] <= r_data[1076];
                
                r_data[1078] <= r_data[1077];
                
                r_data[1079] <= r_data[1078];
                
                r_data[1080] <= r_data[1079];
                
                r_data[1081] <= r_data[1080];
                
                r_data[1082] <= r_data[1081];
                
                r_data[1083] <= r_data[1082];
                
                r_data[1084] <= r_data[1083];
                
                r_data[1085] <= r_data[1084];
                
                r_data[1086] <= r_data[1085];
                
                r_data[1087] <= r_data[1086];
                
                r_data[1088] <= r_data[1087];
                
                r_data[1089] <= r_data[1088];
                
                r_data[1090] <= r_data[1089];
                
                r_data[1091] <= r_data[1090];
                
                r_data[1092] <= r_data[1091];
                
                r_data[1093] <= r_data[1092];
                
                r_data[1094] <= r_data[1093];
                
                r_data[1095] <= r_data[1094];
                
                r_data[1096] <= r_data[1095];
                
                r_data[1097] <= r_data[1096];
                
                r_data[1098] <= r_data[1097];
                
                r_data[1099] <= r_data[1098];
                
                r_data[1100] <= r_data[1099];
                
                r_data[1101] <= r_data[1100];
                
                r_data[1102] <= r_data[1101];
                
                r_data[1103] <= r_data[1102];
                
                r_data[1104] <= r_data[1103];
                
                r_data[1105] <= r_data[1104];
                
                r_data[1106] <= r_data[1105];
                
                r_data[1107] <= r_data[1106];
                
                r_data[1108] <= r_data[1107];
                
                r_data[1109] <= r_data[1108];
                
                r_data[1110] <= r_data[1109];
                
                r_data[1111] <= r_data[1110];
                
                r_data[1112] <= r_data[1111];
                
                r_data[1113] <= r_data[1112];
                
                r_data[1114] <= r_data[1113];
                
                r_data[1115] <= r_data[1114];
                
                r_data[1116] <= r_data[1115];
                
                r_data[1117] <= r_data[1116];
                
                r_data[1118] <= r_data[1117];
                
                r_data[1119] <= r_data[1118];
                
                r_data[1120] <= r_data[1119];
                
                r_data[1121] <= r_data[1120];
                
                r_data[1122] <= r_data[1121];
                
                r_data[1123] <= r_data[1122];
                
                r_data[1124] <= r_data[1123];
                
                r_data[1125] <= r_data[1124];
                
                r_data[1126] <= r_data[1125];
                
                r_data[1127] <= r_data[1126];
                
                r_data[1128] <= r_data[1127];
                
                r_data[1129] <= r_data[1128];
                
                r_data[1130] <= r_data[1129];
                
                r_data[1131] <= r_data[1130];
                
                r_data[1132] <= r_data[1131];
                
                r_data[1133] <= r_data[1132];
                
                r_data[1134] <= r_data[1133];
                
                r_data[1135] <= r_data[1134];
                
                r_data[1136] <= r_data[1135];
                
                r_data[1137] <= r_data[1136];
                
                r_data[1138] <= r_data[1137];
                
                r_data[1139] <= r_data[1138];
                
                r_data[1140] <= r_data[1139];
                
                r_data[1141] <= r_data[1140];
                
                r_data[1142] <= r_data[1141];
                
                r_data[1143] <= r_data[1142];
                
                r_data[1144] <= r_data[1143];
                
                r_data[1145] <= r_data[1144];
                
                r_data[1146] <= r_data[1145];
                
                r_data[1147] <= r_data[1146];
                
                r_data[1148] <= r_data[1147];
                
                r_data[1149] <= r_data[1148];
                
                r_data[1150] <= r_data[1149];
                
                r_data[1151] <= r_data[1150];
                
                r_data[1152] <= r_data[1151];
                
                r_data[1153] <= r_data[1152];
                
                r_data[1154] <= r_data[1153];
                
                r_data[1155] <= r_data[1154];
                
                r_data[1156] <= r_data[1155];
                
                r_data[1157] <= r_data[1156];
                
                r_data[1158] <= r_data[1157];
                
                r_data[1159] <= r_data[1158];
                
                r_data[1160] <= r_data[1159];
                
                r_data[1161] <= r_data[1160];
                
                r_data[1162] <= r_data[1161];
                
                r_data[1163] <= r_data[1162];
                
                r_data[1164] <= r_data[1163];
                
                r_data[1165] <= r_data[1164];
                
                r_data[1166] <= r_data[1165];
                
                r_data[1167] <= r_data[1166];
                
                r_data[1168] <= r_data[1167];
                
                r_data[1169] <= r_data[1168];
                
                r_data[1170] <= r_data[1169];
                
                r_data[1171] <= r_data[1170];
                
                r_data[1172] <= r_data[1171];
                
                r_data[1173] <= r_data[1172];
                
                r_data[1174] <= r_data[1173];
                
                r_data[1175] <= r_data[1174];
                
                r_data[1176] <= r_data[1175];
                
                r_data[1177] <= r_data[1176];
                
                r_data[1178] <= r_data[1177];
                
                r_data[1179] <= r_data[1178];
                
                r_data[1180] <= r_data[1179];
                
                r_data[1181] <= r_data[1180];
                
                r_data[1182] <= r_data[1181];
                
                r_data[1183] <= r_data[1182];
                
                r_data[1184] <= r_data[1183];
                
                r_data[1185] <= r_data[1184];
                
                r_data[1186] <= r_data[1185];
                
                r_data[1187] <= r_data[1186];
                
                r_data[1188] <= r_data[1187];
                
                r_data[1189] <= r_data[1188];
                
                r_data[1190] <= r_data[1189];
                
                r_data[1191] <= r_data[1190];
                
                r_data[1192] <= r_data[1191];
                
                r_data[1193] <= r_data[1192];
                
                r_data[1194] <= r_data[1193];
                
                r_data[1195] <= r_data[1194];
                
                r_data[1196] <= r_data[1195];
                
                r_data[1197] <= r_data[1196];
                
                r_data[1198] <= r_data[1197];
                
                r_data[1199] <= r_data[1198];
                
                r_data[1200] <= r_data[1199];
                
                r_data[1201] <= r_data[1200];
                
                r_data[1202] <= r_data[1201];
                
                r_data[1203] <= r_data[1202];
                
                r_data[1204] <= r_data[1203];
                
                r_data[1205] <= r_data[1204];
                
                r_data[1206] <= r_data[1205];
                
                r_data[1207] <= r_data[1206];
                
                r_data[1208] <= r_data[1207];
                
                r_data[1209] <= r_data[1208];
                
                r_data[1210] <= r_data[1209];
                
                r_data[1211] <= r_data[1210];
                
                r_data[1212] <= r_data[1211];
                
                r_data[1213] <= r_data[1212];
                
                r_data[1214] <= r_data[1213];
                
                r_data[1215] <= r_data[1214];
                
                r_data[1216] <= r_data[1215];
                
                r_data[1217] <= r_data[1216];
                
                r_data[1218] <= r_data[1217];
                
                r_data[1219] <= r_data[1218];
                
                r_data[1220] <= r_data[1219];
                
                r_data[1221] <= r_data[1220];
                
                r_data[1222] <= r_data[1221];
                
                r_data[1223] <= r_data[1222];
                
                r_data[1224] <= r_data[1223];
                
                r_data[1225] <= r_data[1224];
                
                r_data[1226] <= r_data[1225];
                
                r_data[1227] <= r_data[1226];
                
                r_data[1228] <= r_data[1227];
                
                r_data[1229] <= r_data[1228];
                
                r_data[1230] <= r_data[1229];
                
                r_data[1231] <= r_data[1230];
                
                r_data[1232] <= r_data[1231];
                
                r_data[1233] <= r_data[1232];
                
                r_data[1234] <= r_data[1233];
                
                r_data[1235] <= r_data[1234];
                
                r_data[1236] <= r_data[1235];
                
                r_data[1237] <= r_data[1236];
                
                r_data[1238] <= r_data[1237];
                
                r_data[1239] <= r_data[1238];
                
                r_data[1240] <= r_data[1239];
                
                r_data[1241] <= r_data[1240];
                
                r_data[1242] <= r_data[1241];
                
                r_data[1243] <= r_data[1242];
                
                r_data[1244] <= r_data[1243];
                
                r_data[1245] <= r_data[1244];
                
                r_data[1246] <= r_data[1245];
                
                r_data[1247] <= r_data[1246];
                
                r_data[1248] <= r_data[1247];
                
                r_data[1249] <= r_data[1248];
                
                r_data[1250] <= r_data[1249];
                
                r_data[1251] <= r_data[1250];
                
                r_data[1252] <= r_data[1251];
                
                r_data[1253] <= r_data[1252];
                
                r_data[1254] <= r_data[1253];
                
                r_data[1255] <= r_data[1254];
                
                r_data[1256] <= r_data[1255];
                
                r_data[1257] <= r_data[1256];
                
                r_data[1258] <= r_data[1257];
                
                r_data[1259] <= r_data[1258];
                
                r_data[1260] <= r_data[1259];
                
                r_data[1261] <= r_data[1260];
                
                r_data[1262] <= r_data[1261];
                
                r_data[1263] <= r_data[1262];
                
                r_data[1264] <= r_data[1263];
                
                r_data[1265] <= r_data[1264];
                
                r_data[1266] <= r_data[1265];
                
                r_data[1267] <= r_data[1266];
                
                r_data[1268] <= r_data[1267];
                
                r_data[1269] <= r_data[1268];
                
                r_data[1270] <= r_data[1269];
                
                r_data[1271] <= r_data[1270];
                
                r_data[1272] <= r_data[1271];
                
                r_data[1273] <= r_data[1272];
                
                r_data[1274] <= r_data[1273];
                
                r_data[1275] <= r_data[1274];
                
                r_data[1276] <= r_data[1275];
                
                r_data[1277] <= r_data[1276];
                
                r_data[1278] <= r_data[1277];
                
                r_data[1279] <= r_data[1278];
                
                r_data[1280] <= r_data[1279];
                
                r_data[1281] <= r_data[1280];
                
                r_data[1282] <= r_data[1281];
                
                r_data[1283] <= r_data[1282];
                
                r_data[1284] <= r_data[1283];
                
                r_data[1285] <= r_data[1284];
                
                r_data[1286] <= r_data[1285];
                
                r_data[1287] <= r_data[1286];
                
                r_data[1288] <= r_data[1287];
                
                r_data[1289] <= r_data[1288];
                
                r_data[1290] <= r_data[1289];
                
                r_data[1291] <= r_data[1290];
                
                r_data[1292] <= r_data[1291];
                
                r_data[1293] <= r_data[1292];
                
                r_data[1294] <= r_data[1293];
                
                r_data[1295] <= r_data[1294];
                
                r_data[1296] <= r_data[1295];
                
                r_data[1297] <= r_data[1296];
                
                r_data[1298] <= r_data[1297];
                
                r_data[1299] <= r_data[1298];
                
                r_data[1300] <= r_data[1299];
                
                r_data[1301] <= r_data[1300];
                
                r_data[1302] <= r_data[1301];
                
                r_data[1303] <= r_data[1302];
                
                r_data[1304] <= r_data[1303];
                
                r_data[1305] <= r_data[1304];
                
                r_data[1306] <= r_data[1305];
                
                r_data[1307] <= r_data[1306];
                
                r_data[1308] <= r_data[1307];
                
                r_data[1309] <= r_data[1308];
                
                r_data[1310] <= r_data[1309];
                
                r_data[1311] <= r_data[1310];
                
                r_data[1312] <= r_data[1311];
                
                r_data[1313] <= r_data[1312];
                
                r_data[1314] <= r_data[1313];
                
                r_data[1315] <= r_data[1314];
                
                r_data[1316] <= r_data[1315];
                
                r_data[1317] <= r_data[1316];
                
                r_data[1318] <= r_data[1317];
                
                r_data[1319] <= r_data[1318];
                
                r_data[1320] <= r_data[1319];
                
                r_data[1321] <= r_data[1320];
                
                r_data[1322] <= r_data[1321];
                
                r_data[1323] <= r_data[1322];
                
                r_data[1324] <= r_data[1323];
                
                r_data[1325] <= r_data[1324];
                
                r_data[1326] <= r_data[1325];
                
                r_data[1327] <= r_data[1326];
                
                r_data[1328] <= r_data[1327];
                
                r_data[1329] <= r_data[1328];
                
                r_data[1330] <= r_data[1329];
                
                r_data[1331] <= r_data[1330];
                
                r_data[1332] <= r_data[1331];
                
                r_data[1333] <= r_data[1332];
                
                r_data[1334] <= r_data[1333];
                
                r_data[1335] <= r_data[1334];
                
                r_data[1336] <= r_data[1335];
                
                r_data[1337] <= r_data[1336];
                
                r_data[1338] <= r_data[1337];
                
                r_data[1339] <= r_data[1338];
                
                r_data[1340] <= r_data[1339];
                
                r_data[1341] <= r_data[1340];
                
                r_data[1342] <= r_data[1341];
                
                r_data[1343] <= r_data[1342];
                
                r_data[1344] <= r_data[1343];
                
                r_data[1345] <= r_data[1344];
                
                r_data[1346] <= r_data[1345];
                
                r_data[1347] <= r_data[1346];
                
                r_data[1348] <= r_data[1347];
                
                r_data[1349] <= r_data[1348];
                
                r_data[1350] <= r_data[1349];
                
                r_data[1351] <= r_data[1350];
                
                r_data[1352] <= r_data[1351];
                
                r_data[1353] <= r_data[1352];
                
                r_data[1354] <= r_data[1353];
                
                r_data[1355] <= r_data[1354];
                
                r_data[1356] <= r_data[1355];
                
                r_data[1357] <= r_data[1356];
                
                r_data[1358] <= r_data[1357];
                
                r_data[1359] <= r_data[1358];
                
                r_data[1360] <= r_data[1359];
                
                r_data[1361] <= r_data[1360];
                
                r_data[1362] <= r_data[1361];
                
                r_data[1363] <= r_data[1362];
                
                r_data[1364] <= r_data[1363];
                
                r_data[1365] <= r_data[1364];
                
                r_data[1366] <= r_data[1365];
                
                r_data[1367] <= r_data[1366];
                
                r_data[1368] <= r_data[1367];
                
                r_data[1369] <= r_data[1368];
                
                r_data[1370] <= r_data[1369];
                
                r_data[1371] <= r_data[1370];
                
                r_data[1372] <= r_data[1371];
                
                r_data[1373] <= r_data[1372];
                
                r_data[1374] <= r_data[1373];
                
                r_data[1375] <= r_data[1374];
                
                r_data[1376] <= r_data[1375];
                
                r_data[1377] <= r_data[1376];
                
                r_data[1378] <= r_data[1377];
                
                r_data[1379] <= r_data[1378];
                
                r_data[1380] <= r_data[1379];
                
                r_data[1381] <= r_data[1380];
                
                r_data[1382] <= r_data[1381];
                
                r_data[1383] <= r_data[1382];
                
                r_data[1384] <= r_data[1383];
                
                r_data[1385] <= r_data[1384];
                
                r_data[1386] <= r_data[1385];
                
                r_data[1387] <= r_data[1386];
                
                r_data[1388] <= r_data[1387];
                
                r_data[1389] <= r_data[1388];
                
                r_data[1390] <= r_data[1389];
                
                r_data[1391] <= r_data[1390];
                
                r_data[1392] <= r_data[1391];
                
                r_data[1393] <= r_data[1392];
                
                r_data[1394] <= r_data[1393];
                
                r_data[1395] <= r_data[1394];
                
                r_data[1396] <= r_data[1395];
                
                r_data[1397] <= r_data[1396];
                
                r_data[1398] <= r_data[1397];
                
                r_data[1399] <= r_data[1398];
                
                r_data[1400] <= r_data[1399];
                
                r_data[1401] <= r_data[1400];
                
                r_data[1402] <= r_data[1401];
                
                r_data[1403] <= r_data[1402];
                
                r_data[1404] <= r_data[1403];
                
                r_data[1405] <= r_data[1404];
                
                r_data[1406] <= r_data[1405];
                
                r_data[1407] <= r_data[1406];
                
                r_data[1408] <= r_data[1407];
                
                r_data[1409] <= r_data[1408];
                
                r_data[1410] <= r_data[1409];
                
                r_data[1411] <= r_data[1410];
                
                r_data[1412] <= r_data[1411];
                
                r_data[1413] <= r_data[1412];
                
                r_data[1414] <= r_data[1413];
                
                r_data[1415] <= r_data[1414];
                
                r_data[1416] <= r_data[1415];
                
                r_data[1417] <= r_data[1416];
                
                r_data[1418] <= r_data[1417];
                
                r_data[1419] <= r_data[1418];
                
                r_data[1420] <= r_data[1419];
                
                r_data[1421] <= r_data[1420];
                
                r_data[1422] <= r_data[1421];
                
                r_data[1423] <= r_data[1422];
                
                r_data[1424] <= r_data[1423];
                
                r_data[1425] <= r_data[1424];
                
                r_data[1426] <= r_data[1425];
                
                r_data[1427] <= r_data[1426];
                
                r_data[1428] <= r_data[1427];
                
                r_data[1429] <= r_data[1428];
                
                r_data[1430] <= r_data[1429];
                
                r_data[1431] <= r_data[1430];
                
                r_data[1432] <= r_data[1431];
                
                r_data[1433] <= r_data[1432];
                
                r_data[1434] <= r_data[1433];
                
                r_data[1435] <= r_data[1434];
                
                r_data[1436] <= r_data[1435];
                
                r_data[1437] <= r_data[1436];
                
                r_data[1438] <= r_data[1437];
                
                r_data[1439] <= r_data[1438];
                
                r_data[1440] <= r_data[1439];
                
                r_data[1441] <= r_data[1440];
                
                r_data[1442] <= r_data[1441];
                
                r_data[1443] <= r_data[1442];
                
                r_data[1444] <= r_data[1443];
                
                r_data[1445] <= r_data[1444];
                
                r_data[1446] <= r_data[1445];
                
                r_data[1447] <= r_data[1446];
                
                r_data[1448] <= r_data[1447];
                
                r_data[1449] <= r_data[1448];
                
                r_data[1450] <= r_data[1449];
                
                r_data[1451] <= r_data[1450];
                
                r_data[1452] <= r_data[1451];
                
                r_data[1453] <= r_data[1452];
                
                r_data[1454] <= r_data[1453];
                
                r_data[1455] <= r_data[1454];
                
                r_data[1456] <= r_data[1455];
                
                r_data[1457] <= r_data[1456];
                
                r_data[1458] <= r_data[1457];
                
                r_data[1459] <= r_data[1458];
                
                r_data[1460] <= r_data[1459];
                
                r_data[1461] <= r_data[1460];
                
                r_data[1462] <= r_data[1461];
                
                r_data[1463] <= r_data[1462];
                
                r_data[1464] <= r_data[1463];
                
                r_data[1465] <= r_data[1464];
                
                r_data[1466] <= r_data[1465];
                
                r_data[1467] <= r_data[1466];
                
                r_data[1468] <= r_data[1467];
                
                r_data[1469] <= r_data[1468];
                
                r_data[1470] <= r_data[1469];
                
                r_data[1471] <= r_data[1470];
                
                r_data[1472] <= r_data[1471];
                
                r_data[1473] <= r_data[1472];
                
                r_data[1474] <= r_data[1473];
                
                r_data[1475] <= r_data[1474];
                
                r_data[1476] <= r_data[1475];
                
                r_data[1477] <= r_data[1476];
                
                r_data[1478] <= r_data[1477];
                
                r_data[1479] <= r_data[1478];
                
                r_data[1480] <= r_data[1479];
                
                r_data[1481] <= r_data[1480];
                
                r_data[1482] <= r_data[1481];
                
                r_data[1483] <= r_data[1482];
                
                r_data[1484] <= r_data[1483];
                
                r_data[1485] <= r_data[1484];
                
                r_data[1486] <= r_data[1485];
                
                r_data[1487] <= r_data[1486];
                
                r_data[1488] <= r_data[1487];
                
                r_data[1489] <= r_data[1488];
                
                r_data[1490] <= r_data[1489];
                
                r_data[1491] <= r_data[1490];
                
                r_data[1492] <= r_data[1491];
                
                r_data[1493] <= r_data[1492];
                
                r_data[1494] <= r_data[1493];
                
                r_data[1495] <= r_data[1494];
                
                r_data[1496] <= r_data[1495];
                
                r_data[1497] <= r_data[1496];
                
                r_data[1498] <= r_data[1497];
                
                r_data[1499] <= r_data[1498];
                
                r_data[1500] <= r_data[1499];
                
                r_data[1501] <= r_data[1500];
                
                r_data[1502] <= r_data[1501];
                
                r_data[1503] <= r_data[1502];
                
                r_data[1504] <= r_data[1503];
                
                r_data[1505] <= r_data[1504];
                
                r_data[1506] <= r_data[1505];
                
                r_data[1507] <= r_data[1506];
                
                r_data[1508] <= r_data[1507];
                
                r_data[1509] <= r_data[1508];
                
                r_data[1510] <= r_data[1509];
                
                r_data[1511] <= r_data[1510];
                
                r_data[1512] <= r_data[1511];
                
                r_data[1513] <= r_data[1512];
                
                r_data[1514] <= r_data[1513];
                
                r_data[1515] <= r_data[1514];
                
                r_data[1516] <= r_data[1515];
                
                r_data[1517] <= r_data[1516];
                
                r_data[1518] <= r_data[1517];
                
                r_data[1519] <= r_data[1518];
                
                r_data[1520] <= r_data[1519];
                
                r_data[1521] <= r_data[1520];
                
                r_data[1522] <= r_data[1521];
                
                r_data[1523] <= r_data[1522];
                
                r_data[1524] <= r_data[1523];
                
                r_data[1525] <= r_data[1524];
                
                r_data[1526] <= r_data[1525];
                
                r_data[1527] <= r_data[1526];
                
                r_data[1528] <= r_data[1527];
                
                r_data[1529] <= r_data[1528];
                
                r_data[1530] <= r_data[1529];
                
                r_data[1531] <= r_data[1530];
                
                r_data[1532] <= r_data[1531];
                
                r_data[1533] <= r_data[1532];
                
                r_data[1534] <= r_data[1533];
                
                r_data[1535] <= r_data[1534];
                
                r_data[1536] <= r_data[1535];
                
                r_data[1537] <= r_data[1536];
                
                r_data[1538] <= r_data[1537];
                
                r_data[1539] <= r_data[1538];
                
                r_data[1540] <= r_data[1539];
                
                r_data[1541] <= r_data[1540];
                
                r_data[1542] <= r_data[1541];
                
                r_data[1543] <= r_data[1542];
                
                r_data[1544] <= r_data[1543];
                
                r_data[1545] <= r_data[1544];
                
                r_data[1546] <= r_data[1545];
                
                r_data[1547] <= r_data[1546];
                
                r_data[1548] <= r_data[1547];
                
                r_data[1549] <= r_data[1548];
                
                r_data[1550] <= r_data[1549];
                
                r_data[1551] <= r_data[1550];
                
                r_data[1552] <= r_data[1551];
                
                r_data[1553] <= r_data[1552];
                
                r_data[1554] <= r_data[1553];
                
                r_data[1555] <= r_data[1554];
                
                r_data[1556] <= r_data[1555];
                
                r_data[1557] <= r_data[1556];
                
                r_data[1558] <= r_data[1557];
                
                r_data[1559] <= r_data[1558];
                
                r_data[1560] <= r_data[1559];
                
                r_data[1561] <= r_data[1560];
                
                r_data[1562] <= r_data[1561];
                
                r_data[1563] <= r_data[1562];
                
                r_data[1564] <= r_data[1563];
                
                r_data[1565] <= r_data[1564];
                
                r_data[1566] <= r_data[1565];
                
                r_data[1567] <= r_data[1566];
                
                r_data[1568] <= r_data[1567];
                
                r_data[1569] <= r_data[1568];
                
                r_data[1570] <= r_data[1569];
                
                r_data[1571] <= r_data[1570];
                
                r_data[1572] <= r_data[1571];
                
                r_data[1573] <= r_data[1572];
                
                r_data[1574] <= r_data[1573];
                
                r_data[1575] <= r_data[1574];
                
                r_data[1576] <= r_data[1575];
                
                r_data[1577] <= r_data[1576];
                
                r_data[1578] <= r_data[1577];
                
                r_data[1579] <= r_data[1578];
                
                r_data[1580] <= r_data[1579];
                
                r_data[1581] <= r_data[1580];
                
                r_data[1582] <= r_data[1581];
                
                r_data[1583] <= r_data[1582];
                
                r_data[1584] <= r_data[1583];
                
                r_data[1585] <= r_data[1584];
                
                r_data[1586] <= r_data[1585];
                
                r_data[1587] <= r_data[1586];
                
                r_data[1588] <= r_data[1587];
                
                r_data[1589] <= r_data[1588];
                
                r_data[1590] <= r_data[1589];
                
                r_data[1591] <= r_data[1590];
                
                r_data[1592] <= r_data[1591];
                
                r_data[1593] <= r_data[1592];
                
                r_data[1594] <= r_data[1593];
                
                r_data[1595] <= r_data[1594];
                
                r_data[1596] <= r_data[1595];
                
                r_data[1597] <= r_data[1596];
                
                r_data[1598] <= r_data[1597];
                
                r_data[1599] <= r_data[1598];
                
                r_data[1600] <= r_data[1599];
                
                r_data[1601] <= r_data[1600];
                
                r_data[1602] <= r_data[1601];
                
                r_data[1603] <= r_data[1602];
                
                r_data[1604] <= r_data[1603];
                
                r_data[1605] <= r_data[1604];
                
                r_data[1606] <= r_data[1605];
                
                r_data[1607] <= r_data[1606];
                
                r_data[1608] <= r_data[1607];
                
                r_data[1609] <= r_data[1608];
                
                r_data[1610] <= r_data[1609];
                
                r_data[1611] <= r_data[1610];
                
                r_data[1612] <= r_data[1611];
                
                r_data[1613] <= r_data[1612];
                
                r_data[1614] <= r_data[1613];
                
                r_data[1615] <= r_data[1614];
                
                r_data[1616] <= r_data[1615];
                
                r_data[1617] <= r_data[1616];
                
                r_data[1618] <= r_data[1617];
                
                r_data[1619] <= r_data[1618];
                
                r_data[1620] <= r_data[1619];
                
                r_data[1621] <= r_data[1620];
                
                r_data[1622] <= r_data[1621];
                
                r_data[1623] <= r_data[1622];
                
                r_data[1624] <= r_data[1623];
                
                r_data[1625] <= r_data[1624];
                
                r_data[1626] <= r_data[1625];
                
                r_data[1627] <= r_data[1626];
                
                r_data[1628] <= r_data[1627];
                
                r_data[1629] <= r_data[1628];
                
                r_data[1630] <= r_data[1629];
                
                r_data[1631] <= r_data[1630];
                
                r_data[1632] <= r_data[1631];
                
                r_data[1633] <= r_data[1632];
                
                r_data[1634] <= r_data[1633];
                
                r_data[1635] <= r_data[1634];
                
                r_data[1636] <= r_data[1635];
                
                r_data[1637] <= r_data[1636];
                
                r_data[1638] <= r_data[1637];
                
                r_data[1639] <= r_data[1638];
                
                r_data[1640] <= r_data[1639];
                
                r_data[1641] <= r_data[1640];
                
                r_data[1642] <= r_data[1641];
                
                r_data[1643] <= r_data[1642];
                
                r_data[1644] <= r_data[1643];
                
                r_data[1645] <= r_data[1644];
                
                r_data[1646] <= r_data[1645];
                
                r_data[1647] <= r_data[1646];
                
                r_data[1648] <= r_data[1647];
                
                r_data[1649] <= r_data[1648];
                
                r_data[1650] <= r_data[1649];
                
                r_data[1651] <= r_data[1650];
                
                r_data[1652] <= r_data[1651];
                
                r_data[1653] <= r_data[1652];
                
                r_data[1654] <= r_data[1653];
                
                r_data[1655] <= r_data[1654];
                
                r_data[1656] <= r_data[1655];
                
                r_data[1657] <= r_data[1656];
                
                r_data[1658] <= r_data[1657];
                
                r_data[1659] <= r_data[1658];
                
                r_data[1660] <= r_data[1659];
                
                r_data[1661] <= r_data[1660];
                
                r_data[1662] <= r_data[1661];
                
                r_data[1663] <= r_data[1662];
                
                r_data[1664] <= r_data[1663];
                
                r_data[1665] <= r_data[1664];
                
                r_data[1666] <= r_data[1665];
                
                r_data[1667] <= r_data[1666];
                
                r_data[1668] <= r_data[1667];
                
                r_data[1669] <= r_data[1668];
                
                r_data[1670] <= r_data[1669];
                
                r_data[1671] <= r_data[1670];
                
                r_data[1672] <= r_data[1671];
                
                r_data[1673] <= r_data[1672];
                
                r_data[1674] <= r_data[1673];
                
                r_data[1675] <= r_data[1674];
                
                r_data[1676] <= r_data[1675];
                
                r_data[1677] <= r_data[1676];
                
                r_data[1678] <= r_data[1677];
                
                r_data[1679] <= r_data[1678];
                
                r_data[1680] <= r_data[1679];
                
                r_data[1681] <= r_data[1680];
                
                r_data[1682] <= r_data[1681];
                
                r_data[1683] <= r_data[1682];
                
                r_data[1684] <= r_data[1683];
                
                r_data[1685] <= r_data[1684];
                
                r_data[1686] <= r_data[1685];
                
                r_data[1687] <= r_data[1686];
                
                r_data[1688] <= r_data[1687];
                
                r_data[1689] <= r_data[1688];
                
                r_data[1690] <= r_data[1689];
                
                r_data[1691] <= r_data[1690];
                
                r_data[1692] <= r_data[1691];
                
                r_data[1693] <= r_data[1692];
                
                r_data[1694] <= r_data[1693];
                
                r_data[1695] <= r_data[1694];
                
                r_data[1696] <= r_data[1695];
                
                r_data[1697] <= r_data[1696];
                
                r_data[1698] <= r_data[1697];
                
                r_data[1699] <= r_data[1698];
                
                r_data[1700] <= r_data[1699];
                
                r_data[1701] <= r_data[1700];
                
                r_data[1702] <= r_data[1701];
                
                r_data[1703] <= r_data[1702];
                
                r_data[1704] <= r_data[1703];
                
                r_data[1705] <= r_data[1704];
                
                r_data[1706] <= r_data[1705];
                
                r_data[1707] <= r_data[1706];
                
                r_data[1708] <= r_data[1707];
                
                r_data[1709] <= r_data[1708];
                
                r_data[1710] <= r_data[1709];
                
                r_data[1711] <= r_data[1710];
                
                r_data[1712] <= r_data[1711];
                
                r_data[1713] <= r_data[1712];
                
                r_data[1714] <= r_data[1713];
                
                r_data[1715] <= r_data[1714];
                
                r_data[1716] <= r_data[1715];
                
                r_data[1717] <= r_data[1716];
                
                r_data[1718] <= r_data[1717];
                
                r_data[1719] <= r_data[1718];
                
                r_data[1720] <= r_data[1719];
                
                r_data[1721] <= r_data[1720];
                
                r_data[1722] <= r_data[1721];
                
                r_data[1723] <= r_data[1722];
                
                r_data[1724] <= r_data[1723];
                
                r_data[1725] <= r_data[1724];
                
                r_data[1726] <= r_data[1725];
                
                r_data[1727] <= r_data[1726];
                
                r_data[1728] <= r_data[1727];
                
                r_data[1729] <= r_data[1728];
                
                r_data[1730] <= r_data[1729];
                
                r_data[1731] <= r_data[1730];
                
                r_data[1732] <= r_data[1731];
                
                r_data[1733] <= r_data[1732];
                
                r_data[1734] <= r_data[1733];
                
                r_data[1735] <= r_data[1734];
                
                r_data[1736] <= r_data[1735];
                
                r_data[1737] <= r_data[1736];
                
                r_data[1738] <= r_data[1737];
                
                r_data[1739] <= r_data[1738];
                
                r_data[1740] <= r_data[1739];
                
                r_data[1741] <= r_data[1740];
                
                r_data[1742] <= r_data[1741];
                
                r_data[1743] <= r_data[1742];
                
                r_data[1744] <= r_data[1743];
                
                r_data[1745] <= r_data[1744];
                
                r_data[1746] <= r_data[1745];
                
                r_data[1747] <= r_data[1746];
                
                r_data[1748] <= r_data[1747];
                
                r_data[1749] <= r_data[1748];
                
                r_data[1750] <= r_data[1749];
                
                r_data[1751] <= r_data[1750];
                
                r_data[1752] <= r_data[1751];
                
                r_data[1753] <= r_data[1752];
                
                r_data[1754] <= r_data[1753];
                
                r_data[1755] <= r_data[1754];
                
                r_data[1756] <= r_data[1755];
                
                r_data[1757] <= r_data[1756];
                
                r_data[1758] <= r_data[1757];
                
                r_data[1759] <= r_data[1758];
                
                r_data[1760] <= r_data[1759];
                
                r_data[1761] <= r_data[1760];
                
                r_data[1762] <= r_data[1761];
                
                r_data[1763] <= r_data[1762];
                
                r_data[1764] <= r_data[1763];
                
                r_data[1765] <= r_data[1764];
                
                r_data[1766] <= r_data[1765];
                
                r_data[1767] <= r_data[1766];
                
                r_data[1768] <= r_data[1767];
                
                r_data[1769] <= r_data[1768];
                
                r_data[1770] <= r_data[1769];
                
                r_data[1771] <= r_data[1770];
                
                r_data[1772] <= r_data[1771];
                
                r_data[1773] <= r_data[1772];
                
                r_data[1774] <= r_data[1773];
                
                r_data[1775] <= r_data[1774];
                
                r_data[1776] <= r_data[1775];
                
                r_data[1777] <= r_data[1776];
                
                r_data[1778] <= r_data[1777];
                
                r_data[1779] <= r_data[1778];
                
                r_data[1780] <= r_data[1779];
                
                r_data[1781] <= r_data[1780];
                
                r_data[1782] <= r_data[1781];
                
                r_data[1783] <= r_data[1782];
                
                r_data[1784] <= r_data[1783];
                
                r_data[1785] <= r_data[1784];
                
                r_data[1786] <= r_data[1785];
                
                r_data[1787] <= r_data[1786];
                
                r_data[1788] <= r_data[1787];
                
                r_data[1789] <= r_data[1788];
                
                r_data[1790] <= r_data[1789];
                
                r_data[1791] <= r_data[1790];
                
                r_data[1792] <= r_data[1791];
                
                r_data[1793] <= r_data[1792];
                
                r_data[1794] <= r_data[1793];
                
                r_data[1795] <= r_data[1794];
                
                r_data[1796] <= r_data[1795];
                
                r_data[1797] <= r_data[1796];
                
                r_data[1798] <= r_data[1797];
                
                r_data[1799] <= r_data[1798];
                
                r_data[1800] <= r_data[1799];
                
                r_data[1801] <= r_data[1800];
                
                r_data[1802] <= r_data[1801];
                
                r_data[1803] <= r_data[1802];
                
                r_data[1804] <= r_data[1803];
                
                r_data[1805] <= r_data[1804];
                
                r_data[1806] <= r_data[1805];
                
                r_data[1807] <= r_data[1806];
                
                r_data[1808] <= r_data[1807];
                
                r_data[1809] <= r_data[1808];
                
                r_data[1810] <= r_data[1809];
                
                r_data[1811] <= r_data[1810];
                
                r_data[1812] <= r_data[1811];
                
                r_data[1813] <= r_data[1812];
                
                r_data[1814] <= r_data[1813];
                
                r_data[1815] <= r_data[1814];
                
                r_data[1816] <= r_data[1815];
                
                r_data[1817] <= r_data[1816];
                
                r_data[1818] <= r_data[1817];
                
                r_data[1819] <= r_data[1818];
                
                r_data[1820] <= r_data[1819];
                
                r_data[1821] <= r_data[1820];
                
                r_data[1822] <= r_data[1821];
                
                r_data[1823] <= r_data[1822];
                
                r_data[1824] <= r_data[1823];
                
                r_data[1825] <= r_data[1824];
                
                r_data[1826] <= r_data[1825];
                
                r_data[1827] <= r_data[1826];
                
                r_data[1828] <= r_data[1827];
                
                r_data[1829] <= r_data[1828];
                
                r_data[1830] <= r_data[1829];
                
                r_data[1831] <= r_data[1830];
                
                r_data[1832] <= r_data[1831];
                
                r_data[1833] <= r_data[1832];
                
                r_data[1834] <= r_data[1833];
                
                r_data[1835] <= r_data[1834];
                
                r_data[1836] <= r_data[1835];
                
                r_data[1837] <= r_data[1836];
                
                r_data[1838] <= r_data[1837];
                
                r_data[1839] <= r_data[1838];
                
                r_data[1840] <= r_data[1839];
                
                r_data[1841] <= r_data[1840];
                
                r_data[1842] <= r_data[1841];
                
                r_data[1843] <= r_data[1842];
                
                r_data[1844] <= r_data[1843];
                
                r_data[1845] <= r_data[1844];
                
                r_data[1846] <= r_data[1845];
                
                r_data[1847] <= r_data[1846];
                
                r_data[1848] <= r_data[1847];
                
                r_data[1849] <= r_data[1848];
                
                r_data[1850] <= r_data[1849];
                
                r_data[1851] <= r_data[1850];
                
                r_data[1852] <= r_data[1851];
                
                r_data[1853] <= r_data[1852];
                
                r_data[1854] <= r_data[1853];
                
                r_data[1855] <= r_data[1854];
                
                r_data[1856] <= r_data[1855];
                
                r_data[1857] <= r_data[1856];
                
                r_data[1858] <= r_data[1857];
                
                r_data[1859] <= r_data[1858];
                
                r_data[1860] <= r_data[1859];
                
                r_data[1861] <= r_data[1860];
                
                r_data[1862] <= r_data[1861];
                
                r_data[1863] <= r_data[1862];
                
                r_data[1864] <= r_data[1863];
                
                r_data[1865] <= r_data[1864];
                
                r_data[1866] <= r_data[1865];
                
                r_data[1867] <= r_data[1866];
                
                r_data[1868] <= r_data[1867];
                
                r_data[1869] <= r_data[1868];
                
                r_data[1870] <= r_data[1869];
                
                r_data[1871] <= r_data[1870];
                
                r_data[1872] <= r_data[1871];
                
                r_data[1873] <= r_data[1872];
                
                r_data[1874] <= r_data[1873];
                
                r_data[1875] <= r_data[1874];
                
                r_data[1876] <= r_data[1875];
                
                r_data[1877] <= r_data[1876];
                
                r_data[1878] <= r_data[1877];
                
                r_data[1879] <= r_data[1878];
                
                r_data[1880] <= r_data[1879];
                
                r_data[1881] <= r_data[1880];
                
                r_data[1882] <= r_data[1881];
                
                r_data[1883] <= r_data[1882];
                
                r_data[1884] <= r_data[1883];
                
                r_data[1885] <= r_data[1884];
                
                r_data[1886] <= r_data[1885];
                
                r_data[1887] <= r_data[1886];
                
                r_data[1888] <= r_data[1887];
                
                r_data[1889] <= r_data[1888];
                
                r_data[1890] <= r_data[1889];
                
                r_data[1891] <= r_data[1890];
                
                r_data[1892] <= r_data[1891];
                
                r_data[1893] <= r_data[1892];
                
                r_data[1894] <= r_data[1893];
                
                r_data[1895] <= r_data[1894];
                
                r_data[1896] <= r_data[1895];
                
                r_data[1897] <= r_data[1896];
                
                r_data[1898] <= r_data[1897];
                
                r_data[1899] <= r_data[1898];
                
                r_data[1900] <= r_data[1899];
                
                r_data[1901] <= r_data[1900];
                
                r_data[1902] <= r_data[1901];
                
                r_data[1903] <= r_data[1902];
                
                r_data[1904] <= r_data[1903];
                
                r_data[1905] <= r_data[1904];
                
                r_data[1906] <= r_data[1905];
                
                r_data[1907] <= r_data[1906];
                
                r_data[1908] <= r_data[1907];
                
                r_data[1909] <= r_data[1908];
                
                r_data[1910] <= r_data[1909];
                
                r_data[1911] <= r_data[1910];
                
                r_data[1912] <= r_data[1911];
                
                r_data[1913] <= r_data[1912];
                
                r_data[1914] <= r_data[1913];
                
                r_data[1915] <= r_data[1914];
                
                r_data[1916] <= r_data[1915];
                
                r_data[1917] <= r_data[1916];
                
                r_data[1918] <= r_data[1917];
                
                r_data[1919] <= r_data[1918];
                
                r_data[1920] <= r_data[1919];
                
                r_data[1921] <= r_data[1920];
                
                r_data[1922] <= r_data[1921];
                
                r_data[1923] <= r_data[1922];
                
                r_data[1924] <= r_data[1923];
                
                r_data[1925] <= r_data[1924];
                
                r_data[1926] <= r_data[1925];
                
                r_data[1927] <= r_data[1926];
                
                r_data[1928] <= r_data[1927];
                
                r_data[1929] <= r_data[1928];
                
                r_data[1930] <= r_data[1929];
                
                r_data[1931] <= r_data[1930];
                
                r_data[1932] <= r_data[1931];
                
                r_data[1933] <= r_data[1932];
                
                r_data[1934] <= r_data[1933];
                
                r_data[1935] <= r_data[1934];
                
                r_data[1936] <= r_data[1935];
                
                r_data[1937] <= r_data[1936];
                
                r_data[1938] <= r_data[1937];
                
                r_data[1939] <= r_data[1938];
                
                r_data[1940] <= r_data[1939];
                
                r_data[1941] <= r_data[1940];
                
                r_data[1942] <= r_data[1941];
                
                r_data[1943] <= r_data[1942];
                
                r_data[1944] <= r_data[1943];
                
                r_data[1945] <= r_data[1944];
                
                r_data[1946] <= r_data[1945];
                
                r_data[1947] <= r_data[1946];
                
                r_data[1948] <= r_data[1947];
                
                r_data[1949] <= r_data[1948];
                
                r_data[1950] <= r_data[1949];
                
                r_data[1951] <= r_data[1950];
                
                r_data[1952] <= r_data[1951];
                
                r_data[1953] <= r_data[1952];
                
                r_data[1954] <= r_data[1953];
                
                r_data[1955] <= r_data[1954];
                
                r_data[1956] <= r_data[1955];
                
                r_data[1957] <= r_data[1956];
                
                r_data[1958] <= r_data[1957];
                
                r_data[1959] <= r_data[1958];
                
                r_data[1960] <= r_data[1959];
                
                r_data[1961] <= r_data[1960];
                
                r_data[1962] <= r_data[1961];
                
                r_data[1963] <= r_data[1962];
                
                r_data[1964] <= r_data[1963];
                
                r_data[1965] <= r_data[1964];
                
                r_data[1966] <= r_data[1965];
                
                r_data[1967] <= r_data[1966];
                
                r_data[1968] <= r_data[1967];
                
                r_data[1969] <= r_data[1968];
                
                r_data[1970] <= r_data[1969];
                
                r_data[1971] <= r_data[1970];
                
                r_data[1972] <= r_data[1971];
                
                r_data[1973] <= r_data[1972];
                
                r_data[1974] <= r_data[1973];
                
                r_data[1975] <= r_data[1974];
                
                r_data[1976] <= r_data[1975];
                
                r_data[1977] <= r_data[1976];
                
                r_data[1978] <= r_data[1977];
                
                r_data[1979] <= r_data[1978];
                
                r_data[1980] <= r_data[1979];
                
                r_data[1981] <= r_data[1980];
                
                r_data[1982] <= r_data[1981];
                
                r_data[1983] <= r_data[1982];
                
                r_data[1984] <= r_data[1983];
                
                r_data[1985] <= r_data[1984];
                
                r_data[1986] <= r_data[1985];
                
                r_data[1987] <= r_data[1986];
                
                r_data[1988] <= r_data[1987];
                
                r_data[1989] <= r_data[1988];
                
                r_data[1990] <= r_data[1989];
                
                r_data[1991] <= r_data[1990];
                
                r_data[1992] <= r_data[1991];
                
                r_data[1993] <= r_data[1992];
                
                r_data[1994] <= r_data[1993];
                
                r_data[1995] <= r_data[1994];
                
                r_data[1996] <= r_data[1995];
                
                r_data[1997] <= r_data[1996];
                
                r_data[1998] <= r_data[1997];
                
                r_data[1999] <= r_data[1998];
                
                r_data[2000] <= r_data[1999];
                
                r_data[2001] <= r_data[2000];
                
                r_data[2002] <= r_data[2001];
                
                r_data[2003] <= r_data[2002];
                
                r_data[2004] <= r_data[2003];
                
                r_data[2005] <= r_data[2004];
                
                r_data[2006] <= r_data[2005];
                
                r_data[2007] <= r_data[2006];
                
                r_data[2008] <= r_data[2007];
                
                r_data[2009] <= r_data[2008];
                
                r_data[2010] <= r_data[2009];
                
                r_data[2011] <= r_data[2010];
                
                r_data[2012] <= r_data[2011];
                
                r_data[2013] <= r_data[2012];
                
                r_data[2014] <= r_data[2013];
                
                r_data[2015] <= r_data[2014];
                
                r_data[2016] <= r_data[2015];
                
                r_data[2017] <= r_data[2016];
                
                r_data[2018] <= r_data[2017];
                
                r_data[2019] <= r_data[2018];
                
                r_data[2020] <= r_data[2019];
                
                r_data[2021] <= r_data[2020];
                
                r_data[2022] <= r_data[2021];
                
                r_data[2023] <= r_data[2022];
                
                r_data[2024] <= r_data[2023];
                
                r_data[2025] <= r_data[2024];
                
                r_data[2026] <= r_data[2025];
                
                r_data[2027] <= r_data[2026];
                
                r_data[2028] <= r_data[2027];
                
                r_data[2029] <= r_data[2028];
                
                r_data[2030] <= r_data[2029];
                
                r_data[2031] <= r_data[2030];
                
                r_data[2032] <= r_data[2031];
                
                r_data[2033] <= r_data[2032];
                
                r_data[2034] <= r_data[2033];
                
                r_data[2035] <= r_data[2034];
                
                r_data[2036] <= r_data[2035];
                
                r_data[2037] <= r_data[2036];
                
                r_data[2038] <= r_data[2037];
                
                r_data[2039] <= r_data[2038];
                
                r_data[2040] <= r_data[2039];
                
                r_data[2041] <= r_data[2040];
                
                r_data[2042] <= r_data[2041];
                
                r_data[2043] <= r_data[2042];
                
                r_data[2044] <= r_data[2043];
                
                r_data[2045] <= r_data[2044];
                
                r_data[2046] <= r_data[2045];
                
                r_data[2047] <= r_data[2046];
                
                r_data[2048] <= r_data[2047];
                
                r_data[2049] <= r_data[2048];
                
                r_data[2050] <= r_data[2049];
                
                r_data[2051] <= r_data[2050];
                
                r_data[2052] <= r_data[2051];
                
                r_data[2053] <= r_data[2052];
                
                r_data[2054] <= r_data[2053];
                
                r_data[2055] <= r_data[2054];
                
                r_data[2056] <= r_data[2055];
                
                r_data[2057] <= r_data[2056];
                
                r_data[2058] <= r_data[2057];
                
                r_data[2059] <= r_data[2058];
                
                r_data[2060] <= r_data[2059];
                
                r_data[2061] <= r_data[2060];
                
                r_data[2062] <= r_data[2061];
                
                r_data[2063] <= r_data[2062];
                
                r_data[2064] <= r_data[2063];
                
                r_data[2065] <= r_data[2064];
                
                r_data[2066] <= r_data[2065];
                
                r_data[2067] <= r_data[2066];
                
                r_data[2068] <= r_data[2067];
                
                r_data[2069] <= r_data[2068];
                
                r_data[2070] <= r_data[2069];
                
                r_data[2071] <= r_data[2070];
                
                r_data[2072] <= r_data[2071];
                
                r_data[2073] <= r_data[2072];
                
                r_data[2074] <= r_data[2073];
                
                r_data[2075] <= r_data[2074];
                
                r_data[2076] <= r_data[2075];
                
                r_data[2077] <= r_data[2076];
                
                r_data[2078] <= r_data[2077];
                
                r_data[2079] <= r_data[2078];
                
                r_data[2080] <= r_data[2079];
                
                r_data[2081] <= r_data[2080];
                
                r_data[2082] <= r_data[2081];
                
                r_data[2083] <= r_data[2082];
                
                r_data[2084] <= r_data[2083];
                
                r_data[2085] <= r_data[2084];
                
                r_data[2086] <= r_data[2085];
                
                r_data[2087] <= r_data[2086];
                
                r_data[2088] <= r_data[2087];
                
                r_data[2089] <= r_data[2088];
                
                r_data[2090] <= r_data[2089];
                
                r_data[2091] <= r_data[2090];
                
                r_data[2092] <= r_data[2091];
                
                r_data[2093] <= r_data[2092];
                
                r_data[2094] <= r_data[2093];
                
                r_data[2095] <= r_data[2094];
                
                r_data[2096] <= r_data[2095];
                
                r_data[2097] <= r_data[2096];
                
                r_data[2098] <= r_data[2097];
                
                r_data[2099] <= r_data[2098];
                
                r_data[2100] <= r_data[2099];
                
                r_data[2101] <= r_data[2100];
                
                r_data[2102] <= r_data[2101];
                
                r_data[2103] <= r_data[2102];
                
                r_data[2104] <= r_data[2103];
                
                r_data[2105] <= r_data[2104];
                
                r_data[2106] <= r_data[2105];
                
                r_data[2107] <= r_data[2106];
                
                r_data[2108] <= r_data[2107];
                
                r_data[2109] <= r_data[2108];
                
                r_data[2110] <= r_data[2109];
                
                r_data[2111] <= r_data[2110];
                
                r_data[2112] <= r_data[2111];
                
                r_data[2113] <= r_data[2112];
                
                r_data[2114] <= r_data[2113];
                
                r_data[2115] <= r_data[2114];
                
                r_data[2116] <= r_data[2115];
                
                r_data[2117] <= r_data[2116];
                
                r_data[2118] <= r_data[2117];
                
                r_data[2119] <= r_data[2118];
                
                r_data[2120] <= r_data[2119];
                
                r_data[2121] <= r_data[2120];
                
                r_data[2122] <= r_data[2121];
                
                r_data[2123] <= r_data[2122];
                
                r_data[2124] <= r_data[2123];
                
                r_data[2125] <= r_data[2124];
                
                r_data[2126] <= r_data[2125];
                
                r_data[2127] <= r_data[2126];
                
                r_data[2128] <= r_data[2127];
                
                r_data[2129] <= r_data[2128];
                
                r_data[2130] <= r_data[2129];
                
                r_data[2131] <= r_data[2130];
                
                r_data[2132] <= r_data[2131];
                
                r_data[2133] <= r_data[2132];
                
                r_data[2134] <= r_data[2133];
                
                r_data[2135] <= r_data[2134];
                
                r_data[2136] <= r_data[2135];
                
                r_data[2137] <= r_data[2136];
                
                r_data[2138] <= r_data[2137];
                
                r_data[2139] <= r_data[2138];
                
                r_data[2140] <= r_data[2139];
                
                r_data[2141] <= r_data[2140];
                
                r_data[2142] <= r_data[2141];
                
                r_data[2143] <= r_data[2142];
                
                r_data[2144] <= r_data[2143];
                
                r_data[2145] <= r_data[2144];
                
                r_data[2146] <= r_data[2145];
                
                r_data[2147] <= r_data[2146];
                
                r_data[2148] <= r_data[2147];
                
                r_data[2149] <= r_data[2148];
                
                r_data[2150] <= r_data[2149];
                
                r_data[2151] <= r_data[2150];
                
                r_data[2152] <= r_data[2151];
                
                r_data[2153] <= r_data[2152];
                
                r_data[2154] <= r_data[2153];
                
                r_data[2155] <= r_data[2154];
                
                r_data[2156] <= r_data[2155];
                
                r_data[2157] <= r_data[2156];
                
                r_data[2158] <= r_data[2157];
                
                r_data[2159] <= r_data[2158];
                
                r_data[2160] <= r_data[2159];
                
                r_data[2161] <= r_data[2160];
                
                r_data[2162] <= r_data[2161];
                
                r_data[2163] <= r_data[2162];
                
                r_data[2164] <= r_data[2163];
                
                r_data[2165] <= r_data[2164];
                
                r_data[2166] <= r_data[2165];
                
                r_data[2167] <= r_data[2166];
                
                r_data[2168] <= r_data[2167];
                
                r_data[2169] <= r_data[2168];
                
                r_data[2170] <= r_data[2169];
                
                r_data[2171] <= r_data[2170];
                
                r_data[2172] <= r_data[2171];
                
                r_data[2173] <= r_data[2172];
                
                r_data[2174] <= r_data[2173];
                
                r_data[2175] <= r_data[2174];
                
                r_data[2176] <= r_data[2175];
                
                r_data[2177] <= r_data[2176];
                
                r_data[2178] <= r_data[2177];
                
                r_data[2179] <= r_data[2178];
                
                r_data[2180] <= r_data[2179];
                
                r_data[2181] <= r_data[2180];
                
                r_data[2182] <= r_data[2181];
                
                r_data[2183] <= r_data[2182];
                
                r_data[2184] <= r_data[2183];
                
                r_data[2185] <= r_data[2184];
                
                r_data[2186] <= r_data[2185];
                
                r_data[2187] <= r_data[2186];
                
                r_data[2188] <= r_data[2187];
                
                r_data[2189] <= r_data[2188];
                
                r_data[2190] <= r_data[2189];
                
                r_data[2191] <= r_data[2190];
                
                r_data[2192] <= r_data[2191];
                
                r_data[2193] <= r_data[2192];
                
                r_data[2194] <= r_data[2193];
                
                r_data[2195] <= r_data[2194];
                
                r_data[2196] <= r_data[2195];
                
                r_data[2197] <= r_data[2196];
                
                r_data[2198] <= r_data[2197];
                
                r_data[2199] <= r_data[2198];
                
                r_data[2200] <= r_data[2199];
                
                r_data[2201] <= r_data[2200];
                
                r_data[2202] <= r_data[2201];
                
                r_data[2203] <= r_data[2202];
                
                r_data[2204] <= r_data[2203];
                
                r_data[2205] <= r_data[2204];
                
                r_data[2206] <= r_data[2205];
                
                r_data[2207] <= r_data[2206];
                
                r_data[2208] <= r_data[2207];
                
                r_data[2209] <= r_data[2208];
                
                r_data[2210] <= r_data[2209];
                
                r_data[2211] <= r_data[2210];
                
                r_data[2212] <= r_data[2211];
                
                r_data[2213] <= r_data[2212];
                
                r_data[2214] <= r_data[2213];
                
                r_data[2215] <= r_data[2214];
                
                r_data[2216] <= r_data[2215];
                
                r_data[2217] <= r_data[2216];
                
                r_data[2218] <= r_data[2217];
                
                r_data[2219] <= r_data[2218];
                
                r_data[2220] <= r_data[2219];
                
                r_data[2221] <= r_data[2220];
                
                r_data[2222] <= r_data[2221];
                
                r_data[2223] <= r_data[2222];
                
                r_data[2224] <= r_data[2223];
                
                r_data[2225] <= r_data[2224];
                
                r_data[2226] <= r_data[2225];
                
                r_data[2227] <= r_data[2226];
                
                r_data[2228] <= r_data[2227];
                
                r_data[2229] <= r_data[2228];
                
                r_data[2230] <= r_data[2229];
                
                r_data[2231] <= r_data[2230];
                
                r_data[2232] <= r_data[2231];
                
                r_data[2233] <= r_data[2232];
                
                r_data[2234] <= r_data[2233];
                
                r_data[2235] <= r_data[2234];
                
                r_data[2236] <= r_data[2235];
                
                r_data[2237] <= r_data[2236];
                
                r_data[2238] <= r_data[2237];
                
                r_data[2239] <= r_data[2238];
                
                r_data[2240] <= r_data[2239];
                
                r_data[2241] <= r_data[2240];
                
                r_data[2242] <= r_data[2241];
                
                r_data[2243] <= r_data[2242];
                
                r_data[2244] <= r_data[2243];
                
                r_data[2245] <= r_data[2244];
                
                r_data[2246] <= r_data[2245];
                
                r_data[2247] <= r_data[2246];
                
                r_data[2248] <= r_data[2247];
                
                r_data[2249] <= r_data[2248];
                
                r_data[2250] <= r_data[2249];
                
                r_data[2251] <= r_data[2250];
                
                r_data[2252] <= r_data[2251];
                
                r_data[2253] <= r_data[2252];
                
                r_data[2254] <= r_data[2253];
                
                r_data[2255] <= r_data[2254];
                
                r_data[2256] <= r_data[2255];
                
                r_data[2257] <= r_data[2256];
                
                r_data[2258] <= r_data[2257];
                
                r_data[2259] <= r_data[2258];
                
                r_data[2260] <= r_data[2259];
                
                r_data[2261] <= r_data[2260];
                
                r_data[2262] <= r_data[2261];
                
                r_data[2263] <= r_data[2262];
                
                r_data[2264] <= r_data[2263];
                
                r_data[2265] <= r_data[2264];
                
                r_data[2266] <= r_data[2265];
                
                r_data[2267] <= r_data[2266];
                
                r_data[2268] <= r_data[2267];
                
                r_data[2269] <= r_data[2268];
                
                r_data[2270] <= r_data[2269];
                
                r_data[2271] <= r_data[2270];
                
                r_data[2272] <= r_data[2271];
                
                r_data[2273] <= r_data[2272];
                
                r_data[2274] <= r_data[2273];
                
                r_data[2275] <= r_data[2274];
                
                r_data[2276] <= r_data[2275];
                
                r_data[2277] <= r_data[2276];
                
                r_data[2278] <= r_data[2277];
                
                r_data[2279] <= r_data[2278];
                
                r_data[2280] <= r_data[2279];
                
                r_data[2281] <= r_data[2280];
                
                r_data[2282] <= r_data[2281];
                
                r_data[2283] <= r_data[2282];
                
                r_data[2284] <= r_data[2283];
                
                r_data[2285] <= r_data[2284];
                
                r_data[2286] <= r_data[2285];
                
                r_data[2287] <= r_data[2286];
                
                r_data[2288] <= r_data[2287];
                
                r_data[2289] <= r_data[2288];
                
                r_data[2290] <= r_data[2289];
                
                r_data[2291] <= r_data[2290];
                
                r_data[2292] <= r_data[2291];
                
                r_data[2293] <= r_data[2292];
                
                r_data[2294] <= r_data[2293];
                
                r_data[2295] <= r_data[2294];
                
                r_data[2296] <= r_data[2295];
                
                r_data[2297] <= r_data[2296];
                
                r_data[2298] <= r_data[2297];
                
                r_data[2299] <= r_data[2298];
                
                r_data[2300] <= r_data[2299];
                
                r_data[2301] <= r_data[2300];
                
                r_data[2302] <= r_data[2301];
                
                r_data[2303] <= r_data[2302];
                
                r_data[2304] <= r_data[2303];
                
                r_data[2305] <= r_data[2304];
                
                r_data[2306] <= r_data[2305];
                
                r_data[2307] <= r_data[2306];
                
                r_data[2308] <= r_data[2307];
                
                r_data[2309] <= r_data[2308];
                
                r_data[2310] <= r_data[2309];
                
                r_data[2311] <= r_data[2310];
                
                r_data[2312] <= r_data[2311];
                
                r_data[2313] <= r_data[2312];
                
                r_data[2314] <= r_data[2313];
                
                r_data[2315] <= r_data[2314];
                
                r_data[2316] <= r_data[2315];
                
                r_data[2317] <= r_data[2316];
                
                r_data[2318] <= r_data[2317];
                
                r_data[2319] <= r_data[2318];
                
                r_data[2320] <= r_data[2319];
                
                r_data[2321] <= r_data[2320];
                
                r_data[2322] <= r_data[2321];
                
                r_data[2323] <= r_data[2322];
                
                r_data[2324] <= r_data[2323];
                
                r_data[2325] <= r_data[2324];
                
                r_data[2326] <= r_data[2325];
                
                r_data[2327] <= r_data[2326];
                
                r_data[2328] <= r_data[2327];
                
                r_data[2329] <= r_data[2328];
                
                r_data[2330] <= r_data[2329];
                
                r_data[2331] <= r_data[2330];
                
                r_data[2332] <= r_data[2331];
                
                r_data[2333] <= r_data[2332];
                
                r_data[2334] <= r_data[2333];
                
                r_data[2335] <= r_data[2334];
                
                r_data[2336] <= r_data[2335];
                
                r_data[2337] <= r_data[2336];
                
                r_data[2338] <= r_data[2337];
                
                r_data[2339] <= r_data[2338];
                
                r_data[2340] <= r_data[2339];
                
                r_data[2341] <= r_data[2340];
                
                r_data[2342] <= r_data[2341];
                
                r_data[2343] <= r_data[2342];
                
                r_data[2344] <= r_data[2343];
                
                r_data[2345] <= r_data[2344];
                
                r_data[2346] <= r_data[2345];
                
                r_data[2347] <= r_data[2346];
                
                r_data[2348] <= r_data[2347];
                
                r_data[2349] <= r_data[2348];
                
                r_data[2350] <= r_data[2349];
                
                r_data[2351] <= r_data[2350];
                
                r_data[2352] <= r_data[2351];
                
                r_data[2353] <= r_data[2352];
                
                r_data[2354] <= r_data[2353];
                
                r_data[2355] <= r_data[2354];
                
                r_data[2356] <= r_data[2355];
                
                r_data[2357] <= r_data[2356];
                
                r_data[2358] <= r_data[2357];
                
                r_data[2359] <= r_data[2358];
                
                r_data[2360] <= r_data[2359];
                
                r_data[2361] <= r_data[2360];
                
                r_data[2362] <= r_data[2361];
                
                r_data[2363] <= r_data[2362];
                
                r_data[2364] <= r_data[2363];
                
                r_data[2365] <= r_data[2364];
                
                r_data[2366] <= r_data[2365];
                
                r_data[2367] <= r_data[2366];
                
                r_data[2368] <= r_data[2367];
                
                r_data[2369] <= r_data[2368];
                
                r_data[2370] <= r_data[2369];
                
                r_data[2371] <= r_data[2370];
                
                r_data[2372] <= r_data[2371];
                
                r_data[2373] <= r_data[2372];
                
                r_data[2374] <= r_data[2373];
                
                r_data[2375] <= r_data[2374];
                
                r_data[2376] <= r_data[2375];
                
                r_data[2377] <= r_data[2376];
                
                r_data[2378] <= r_data[2377];
                
                r_data[2379] <= r_data[2378];
                
                r_data[2380] <= r_data[2379];
                
                r_data[2381] <= r_data[2380];
                
                r_data[2382] <= r_data[2381];
                
                r_data[2383] <= r_data[2382];
                
                r_data[2384] <= r_data[2383];
                
                r_data[2385] <= r_data[2384];
                
                r_data[2386] <= r_data[2385];
                
                r_data[2387] <= r_data[2386];
                
                r_data[2388] <= r_data[2387];
                
                r_data[2389] <= r_data[2388];
                
                r_data[2390] <= r_data[2389];
                
                r_data[2391] <= r_data[2390];
                
                r_data[2392] <= r_data[2391];
                
                r_data[2393] <= r_data[2392];
                
                r_data[2394] <= r_data[2393];
                
                r_data[2395] <= r_data[2394];
                
                r_data[2396] <= r_data[2395];
                
                r_data[2397] <= r_data[2396];
                
                r_data[2398] <= r_data[2397];
                
                r_data[2399] <= r_data[2398];
                
                r_data[2400] <= r_data[2399];
                
                r_data[2401] <= r_data[2400];
                
                r_data[2402] <= r_data[2401];
                
                r_data[2403] <= r_data[2402];
                
                r_data[2404] <= r_data[2403];
                
                r_data[2405] <= r_data[2404];
                
                r_data[2406] <= r_data[2405];
                
                r_data[2407] <= r_data[2406];
                
                r_data[2408] <= r_data[2407];
                
                r_data[2409] <= r_data[2408];
                
                r_data[2410] <= r_data[2409];
                
                r_data[2411] <= r_data[2410];
                
                r_data[2412] <= r_data[2411];
                
                r_data[2413] <= r_data[2412];
                
                r_data[2414] <= r_data[2413];
                
                r_data[2415] <= r_data[2414];
                
                r_data[2416] <= r_data[2415];
                
                r_data[2417] <= r_data[2416];
                
                r_data[2418] <= r_data[2417];
                
                r_data[2419] <= r_data[2418];
                
                r_data[2420] <= r_data[2419];
                
                r_data[2421] <= r_data[2420];
                
                r_data[2422] <= r_data[2421];
                
                r_data[2423] <= r_data[2422];
                
                r_data[2424] <= r_data[2423];
                
                r_data[2425] <= r_data[2424];
                
                r_data[2426] <= r_data[2425];
                
                r_data[2427] <= r_data[2426];
                
                r_data[2428] <= r_data[2427];
                
                r_data[2429] <= r_data[2428];
                
                r_data[2430] <= r_data[2429];
                
                r_data[2431] <= r_data[2430];
                
                r_data[2432] <= r_data[2431];
                
                r_data[2433] <= r_data[2432];
                
                r_data[2434] <= r_data[2433];
                
                r_data[2435] <= r_data[2434];
                
                r_data[2436] <= r_data[2435];
                
                r_data[2437] <= r_data[2436];
                
                r_data[2438] <= r_data[2437];
                
                r_data[2439] <= r_data[2438];
                
                r_data[2440] <= r_data[2439];
                
                r_data[2441] <= r_data[2440];
                
                r_data[2442] <= r_data[2441];
                
                r_data[2443] <= r_data[2442];
                
                r_data[2444] <= r_data[2443];
                
                r_data[2445] <= r_data[2444];
                
                r_data[2446] <= r_data[2445];
                
                r_data[2447] <= r_data[2446];
                
                r_data[2448] <= r_data[2447];
                
                r_data[2449] <= r_data[2448];
                
                r_data[2450] <= r_data[2449];
                
                r_data[2451] <= r_data[2450];
                
                r_data[2452] <= r_data[2451];
                
                r_data[2453] <= r_data[2452];
                
                r_data[2454] <= r_data[2453];
                
                r_data[2455] <= r_data[2454];
                
                r_data[2456] <= r_data[2455];
                
                r_data[2457] <= r_data[2456];
                
                r_data[2458] <= r_data[2457];
                
                r_data[2459] <= r_data[2458];
                
                r_data[2460] <= r_data[2459];
                
                r_data[2461] <= r_data[2460];
                
                r_data[2462] <= r_data[2461];
                
                r_data[2463] <= r_data[2462];
                
                r_data[2464] <= r_data[2463];
                
                r_data[2465] <= r_data[2464];
                
                r_data[2466] <= r_data[2465];
                
                r_data[2467] <= r_data[2466];
                
                r_data[2468] <= r_data[2467];
                
                r_data[2469] <= r_data[2468];
                
                r_data[2470] <= r_data[2469];
                
                r_data[2471] <= r_data[2470];
                
                r_data[2472] <= r_data[2471];
                
                r_data[2473] <= r_data[2472];
                
                r_data[2474] <= r_data[2473];
                
                r_data[2475] <= r_data[2474];
                
                r_data[2476] <= r_data[2475];
                
                r_data[2477] <= r_data[2476];
                
                r_data[2478] <= r_data[2477];
                
                r_data[2479] <= r_data[2478];
                
                r_data[2480] <= r_data[2479];
                
                r_data[2481] <= r_data[2480];
                
                r_data[2482] <= r_data[2481];
                
                r_data[2483] <= r_data[2482];
                
                r_data[2484] <= r_data[2483];
                
                r_data[2485] <= r_data[2484];
                
                r_data[2486] <= r_data[2485];
                
                r_data[2487] <= r_data[2486];
                
                r_data[2488] <= r_data[2487];
                
                r_data[2489] <= r_data[2488];
                
                r_data[2490] <= r_data[2489];
                
                r_data[2491] <= r_data[2490];
                
                r_data[2492] <= r_data[2491];
                
                r_data[2493] <= r_data[2492];
                
                r_data[2494] <= r_data[2493];
                
                r_data[2495] <= r_data[2494];
                
                r_data[2496] <= r_data[2495];
                
                r_data[2497] <= r_data[2496];
                
                r_data[2498] <= r_data[2497];
                
                r_data[2499] <= r_data[2498];
                
                r_data[2500] <= r_data[2499];
                
                r_data[2501] <= r_data[2500];
                
                r_data[2502] <= r_data[2501];
                
                r_data[2503] <= r_data[2502];
                
                r_data[2504] <= r_data[2503];
                
                r_data[2505] <= r_data[2504];
                
                r_data[2506] <= r_data[2505];
                
                r_data[2507] <= r_data[2506];
                
                r_data[2508] <= r_data[2507];
                
                r_data[2509] <= r_data[2508];
                
                r_data[2510] <= r_data[2509];
                
                r_data[2511] <= r_data[2510];
                
                r_data[2512] <= r_data[2511];
                
                r_data[2513] <= r_data[2512];
                
                r_data[2514] <= r_data[2513];
                
                r_data[2515] <= r_data[2514];
                
                r_data[2516] <= r_data[2515];
                
                r_data[2517] <= r_data[2516];
                
                r_data[2518] <= r_data[2517];
                
                r_data[2519] <= r_data[2518];
                
                r_data[2520] <= r_data[2519];
                
                r_data[2521] <= r_data[2520];
                
                r_data[2522] <= r_data[2521];
                
                r_data[2523] <= r_data[2522];
                
                r_data[2524] <= r_data[2523];
                
                r_data[2525] <= r_data[2524];
                
                r_data[2526] <= r_data[2525];
                
                r_data[2527] <= r_data[2526];
                
                r_data[2528] <= r_data[2527];
                
                r_data[2529] <= r_data[2528];
                
                r_data[2530] <= r_data[2529];
                
                r_data[2531] <= r_data[2530];
                
                r_data[2532] <= r_data[2531];
                
                r_data[2533] <= r_data[2532];
                
                r_data[2534] <= r_data[2533];
                
                r_data[2535] <= r_data[2534];
                
                r_data[2536] <= r_data[2535];
                
                r_data[2537] <= r_data[2536];
                
                r_data[2538] <= r_data[2537];
                
                r_data[2539] <= r_data[2538];
                
                r_data[2540] <= r_data[2539];
                
                r_data[2541] <= r_data[2540];
                
                r_data[2542] <= r_data[2541];
                
                r_data[2543] <= r_data[2542];
                
                r_data[2544] <= r_data[2543];
                
                r_data[2545] <= r_data[2544];
                
                r_data[2546] <= r_data[2545];
                
                r_data[2547] <= r_data[2546];
                
                r_data[2548] <= r_data[2547];
                
                r_data[2549] <= r_data[2548];
                
                r_data[2550] <= r_data[2549];
                
                r_data[2551] <= r_data[2550];
                
                r_data[2552] <= r_data[2551];
                
                r_data[2553] <= r_data[2552];
                
                r_data[2554] <= r_data[2553];
                
                r_data[2555] <= r_data[2554];
                
                r_data[2556] <= r_data[2555];
                
                r_data[2557] <= r_data[2556];
                
                r_data[2558] <= r_data[2557];
                
                r_data[2559] <= r_data[2558];
                
                r_data[2560] <= r_data[2559];
                
                r_data[2561] <= r_data[2560];
                
                r_data[2562] <= r_data[2561];
                
                r_data[2563] <= r_data[2562];
                
                r_data[2564] <= r_data[2563];
                
                r_data[2565] <= r_data[2564];
                
                r_data[2566] <= r_data[2565];
                
                r_data[2567] <= r_data[2566];
                
                r_data[2568] <= r_data[2567];
                
                r_data[2569] <= r_data[2568];
                
                r_data[2570] <= r_data[2569];
                
                r_data[2571] <= r_data[2570];
                
                r_data[2572] <= r_data[2571];
                
                r_data[2573] <= r_data[2572];
                
                r_data[2574] <= r_data[2573];
                
                r_data[2575] <= r_data[2574];
                
                r_data[2576] <= r_data[2575];
                
                r_data[2577] <= r_data[2576];
                
                r_data[2578] <= r_data[2577];
                
                r_data[2579] <= r_data[2578];
                
                r_data[2580] <= r_data[2579];
                
                r_data[2581] <= r_data[2580];
                
                r_data[2582] <= r_data[2581];
                
                r_data[2583] <= r_data[2582];
                
                r_data[2584] <= r_data[2583];
                
                r_data[2585] <= r_data[2584];
                
                r_data[2586] <= r_data[2585];
                
                r_data[2587] <= r_data[2586];
                
                r_data[2588] <= r_data[2587];
                
                r_data[2589] <= r_data[2588];
                
                r_data[2590] <= r_data[2589];
                
                r_data[2591] <= r_data[2590];
                
                r_data[2592] <= r_data[2591];
                
                r_data[2593] <= r_data[2592];
                
                r_data[2594] <= r_data[2593];
                
                r_data[2595] <= r_data[2594];
                
                r_data[2596] <= r_data[2595];
                
                r_data[2597] <= r_data[2596];
                
                r_data[2598] <= r_data[2597];
                
                r_data[2599] <= r_data[2598];
                
                r_data[2600] <= r_data[2599];
                
                r_data[2601] <= r_data[2600];
                
                r_data[2602] <= r_data[2601];
                
                r_data[2603] <= r_data[2602];
                
                r_data[2604] <= r_data[2603];
                
                r_data[2605] <= r_data[2604];
                
                r_data[2606] <= r_data[2605];
                
                r_data[2607] <= r_data[2606];
                
                r_data[2608] <= r_data[2607];
                
                r_data[2609] <= r_data[2608];
                
                r_data[2610] <= r_data[2609];
                
                r_data[2611] <= r_data[2610];
                
                r_data[2612] <= r_data[2611];
                
                r_data[2613] <= r_data[2612];
                
                r_data[2614] <= r_data[2613];
                
                r_data[2615] <= r_data[2614];
                
                r_data[2616] <= r_data[2615];
                
                r_data[2617] <= r_data[2616];
                
                r_data[2618] <= r_data[2617];
                
                r_data[2619] <= r_data[2618];
                
                r_data[2620] <= r_data[2619];
                
                r_data[2621] <= r_data[2620];
                
                r_data[2622] <= r_data[2621];
                
                r_data[2623] <= r_data[2622];
                
                r_data[2624] <= r_data[2623];
                
                r_data[2625] <= r_data[2624];
                
                r_data[2626] <= r_data[2625];
                
                r_data[2627] <= r_data[2626];
                
                r_data[2628] <= r_data[2627];
                
                r_data[2629] <= r_data[2628];
                
                r_data[2630] <= r_data[2629];
                
                r_data[2631] <= r_data[2630];
                
                r_data[2632] <= r_data[2631];
                
                r_data[2633] <= r_data[2632];
                
                r_data[2634] <= r_data[2633];
                
                r_data[2635] <= r_data[2634];
                
                r_data[2636] <= r_data[2635];
                
                r_data[2637] <= r_data[2636];
                
                r_data[2638] <= r_data[2637];
                
                r_data[2639] <= r_data[2638];
                
                r_data[2640] <= r_data[2639];
                
                r_data[2641] <= r_data[2640];
                
                r_data[2642] <= r_data[2641];
                
                r_data[2643] <= r_data[2642];
                
                r_data[2644] <= r_data[2643];
                
                r_data[2645] <= r_data[2644];
                
                r_data[2646] <= r_data[2645];
                
                r_data[2647] <= r_data[2646];
                
                r_data[2648] <= r_data[2647];
                
                r_data[2649] <= r_data[2648];
                
                r_data[2650] <= r_data[2649];
                
                r_data[2651] <= r_data[2650];
                
                r_data[2652] <= r_data[2651];
                
                r_data[2653] <= r_data[2652];
                
                r_data[2654] <= r_data[2653];
                
                r_data[2655] <= r_data[2654];
                
                r_data[2656] <= r_data[2655];
                
                r_data[2657] <= r_data[2656];
                
                r_data[2658] <= r_data[2657];
                
                r_data[2659] <= r_data[2658];
                
                r_data[2660] <= r_data[2659];
                
                r_data[2661] <= r_data[2660];
                
                r_data[2662] <= r_data[2661];
                
                r_data[2663] <= r_data[2662];
                
                r_data[2664] <= r_data[2663];
                
                r_data[2665] <= r_data[2664];
                
                r_data[2666] <= r_data[2665];
                
                r_data[2667] <= r_data[2666];
                
                r_data[2668] <= r_data[2667];
                
                r_data[2669] <= r_data[2668];
                
                r_data[2670] <= r_data[2669];
                
                r_data[2671] <= r_data[2670];
                
                r_data[2672] <= r_data[2671];
                
                r_data[2673] <= r_data[2672];
                
                r_data[2674] <= r_data[2673];
                
                r_data[2675] <= r_data[2674];
                
                r_data[2676] <= r_data[2675];
                
                r_data[2677] <= r_data[2676];
                
                r_data[2678] <= r_data[2677];
                
                r_data[2679] <= r_data[2678];
                
                r_data[2680] <= r_data[2679];
                
                r_data[2681] <= r_data[2680];
                
                r_data[2682] <= r_data[2681];
                
                r_data[2683] <= r_data[2682];
                
                r_data[2684] <= r_data[2683];
                
                r_data[2685] <= r_data[2684];
                
                r_data[2686] <= r_data[2685];
                
                r_data[2687] <= r_data[2686];
                
                r_data[2688] <= r_data[2687];
                
                r_data[2689] <= r_data[2688];
                
                r_data[2690] <= r_data[2689];
                
                r_data[2691] <= r_data[2690];
                
                r_data[2692] <= r_data[2691];
                
                r_data[2693] <= r_data[2692];
                
                r_data[2694] <= r_data[2693];
                
                r_data[2695] <= r_data[2694];
                
                r_data[2696] <= r_data[2695];
                
                r_data[2697] <= r_data[2696];
                
                r_data[2698] <= r_data[2697];
                
                r_data[2699] <= r_data[2698];
                
                r_data[2700] <= r_data[2699];
                
                r_data[2701] <= r_data[2700];
                
                r_data[2702] <= r_data[2701];
                
                r_data[2703] <= r_data[2702];
                
                r_data[2704] <= r_data[2703];
                
                r_data[2705] <= r_data[2704];
                
                r_data[2706] <= r_data[2705];
                
                r_data[2707] <= r_data[2706];
                
                r_data[2708] <= r_data[2707];
                
                r_data[2709] <= r_data[2708];
                
                r_data[2710] <= r_data[2709];
                
                r_data[2711] <= r_data[2710];
                
                r_data[2712] <= r_data[2711];
                
                r_data[2713] <= r_data[2712];
                
                r_data[2714] <= r_data[2713];
                
                r_data[2715] <= r_data[2714];
                
                r_data[2716] <= r_data[2715];
                
                r_data[2717] <= r_data[2716];
                
                r_data[2718] <= r_data[2717];
                
                r_data[2719] <= r_data[2718];
                
                r_data[2720] <= r_data[2719];
                
                r_data[2721] <= r_data[2720];
                
                r_data[2722] <= r_data[2721];
                
                r_data[2723] <= r_data[2722];
                
                r_data[2724] <= r_data[2723];
                
                r_data[2725] <= r_data[2724];
                
                r_data[2726] <= r_data[2725];
                
                r_data[2727] <= r_data[2726];
                
                r_data[2728] <= r_data[2727];
                
                r_data[2729] <= r_data[2728];
                
                r_data[2730] <= r_data[2729];
                
                r_data[2731] <= r_data[2730];
                
                r_data[2732] <= r_data[2731];
                
                r_data[2733] <= r_data[2732];
                
                r_data[2734] <= r_data[2733];
                
                r_data[2735] <= r_data[2734];
                
                r_data[2736] <= r_data[2735];
                
                r_data[2737] <= r_data[2736];
                
                r_data[2738] <= r_data[2737];
                
                r_data[2739] <= r_data[2738];
                
                r_data[2740] <= r_data[2739];
                
                r_data[2741] <= r_data[2740];
                
                r_data[2742] <= r_data[2741];
                
                r_data[2743] <= r_data[2742];
                
                r_data[2744] <= r_data[2743];
                
                r_data[2745] <= r_data[2744];
                
                r_data[2746] <= r_data[2745];
                
                r_data[2747] <= r_data[2746];
                
                r_data[2748] <= r_data[2747];
                
                r_data[2749] <= r_data[2748];
                
                r_data[2750] <= r_data[2749];
                
                r_data[2751] <= r_data[2750];
                
                r_data[2752] <= r_data[2751];
                
                r_data[2753] <= r_data[2752];
                
                r_data[2754] <= r_data[2753];
                
                r_data[2755] <= r_data[2754];
                
                r_data[2756] <= r_data[2755];
                
                r_data[2757] <= r_data[2756];
                
                r_data[2758] <= r_data[2757];
                
                r_data[2759] <= r_data[2758];
                
                r_data[2760] <= r_data[2759];
                
                r_data[2761] <= r_data[2760];
                
                r_data[2762] <= r_data[2761];
                
                r_data[2763] <= r_data[2762];
                
                r_data[2764] <= r_data[2763];
                
                r_data[2765] <= r_data[2764];
                
                r_data[2766] <= r_data[2765];
                
                r_data[2767] <= r_data[2766];
                
                r_data[2768] <= r_data[2767];
                
                r_data[2769] <= r_data[2768];
                
                r_data[2770] <= r_data[2769];
                
                r_data[2771] <= r_data[2770];
                
                r_data[2772] <= r_data[2771];
                
                r_data[2773] <= r_data[2772];
                
                r_data[2774] <= r_data[2773];
                
                r_data[2775] <= r_data[2774];
                
                r_data[2776] <= r_data[2775];
                
                r_data[2777] <= r_data[2776];
                
                r_data[2778] <= r_data[2777];
                
                r_data[2779] <= r_data[2778];
                
                r_data[2780] <= r_data[2779];
                
                r_data[2781] <= r_data[2780];
                
                r_data[2782] <= r_data[2781];
                
                r_data[2783] <= r_data[2782];
                
                r_data[2784] <= r_data[2783];
                
                r_data[2785] <= r_data[2784];
                
                r_data[2786] <= r_data[2785];
                
                r_data[2787] <= r_data[2786];
                
                r_data[2788] <= r_data[2787];
                
                r_data[2789] <= r_data[2788];
                
                r_data[2790] <= r_data[2789];
                
                r_data[2791] <= r_data[2790];
                
                r_data[2792] <= r_data[2791];
                
                r_data[2793] <= r_data[2792];
                
                r_data[2794] <= r_data[2793];
                
                r_data[2795] <= r_data[2794];
                
                r_data[2796] <= r_data[2795];
                
                r_data[2797] <= r_data[2796];
                
                r_data[2798] <= r_data[2797];
                
                r_data[2799] <= r_data[2798];
                
                r_data[2800] <= r_data[2799];
                
                r_data[2801] <= r_data[2800];
                
                r_data[2802] <= r_data[2801];
                
                r_data[2803] <= r_data[2802];
                
                r_data[2804] <= r_data[2803];
                
                r_data[2805] <= r_data[2804];
                
                r_data[2806] <= r_data[2805];
                
                r_data[2807] <= r_data[2806];
                
                r_data[2808] <= r_data[2807];
                
                r_data[2809] <= r_data[2808];
                
                r_data[2810] <= r_data[2809];
                
                r_data[2811] <= r_data[2810];
                
                r_data[2812] <= r_data[2811];
                
                r_data[2813] <= r_data[2812];
                
                r_data[2814] <= r_data[2813];
                
                r_data[2815] <= r_data[2814];
                
                r_data[2816] <= r_data[2815];
                
                r_data[2817] <= r_data[2816];
                
                r_data[2818] <= r_data[2817];
                
                r_data[2819] <= r_data[2818];
                
                r_data[2820] <= r_data[2819];
                
                r_data[2821] <= r_data[2820];
                
                r_data[2822] <= r_data[2821];
                
                r_data[2823] <= r_data[2822];
                
                r_data[2824] <= r_data[2823];
                
                r_data[2825] <= r_data[2824];
                
                r_data[2826] <= r_data[2825];
                
                r_data[2827] <= r_data[2826];
                
                r_data[2828] <= r_data[2827];
                
                r_data[2829] <= r_data[2828];
                
                r_data[2830] <= r_data[2829];
                
                r_data[2831] <= r_data[2830];
                
                r_data[2832] <= r_data[2831];
                
                r_data[2833] <= r_data[2832];
                
                r_data[2834] <= r_data[2833];
                
                r_data[2835] <= r_data[2834];
                
                r_data[2836] <= r_data[2835];
                
                r_data[2837] <= r_data[2836];
                
                r_data[2838] <= r_data[2837];
                
                r_data[2839] <= r_data[2838];
                
                r_data[2840] <= r_data[2839];
                
                r_data[2841] <= r_data[2840];
                
                r_data[2842] <= r_data[2841];
                
                r_data[2843] <= r_data[2842];
                
                r_data[2844] <= r_data[2843];
                
                r_data[2845] <= r_data[2844];
                
                r_data[2846] <= r_data[2845];
                
                r_data[2847] <= r_data[2846];
                
                r_data[2848] <= r_data[2847];
                
                r_data[2849] <= r_data[2848];
                
                r_data[2850] <= r_data[2849];
                
                r_data[2851] <= r_data[2850];
                
                r_data[2852] <= r_data[2851];
                
                r_data[2853] <= r_data[2852];
                
                r_data[2854] <= r_data[2853];
                
                r_data[2855] <= r_data[2854];
                
                r_data[2856] <= r_data[2855];
                
                r_data[2857] <= r_data[2856];
                
                r_data[2858] <= r_data[2857];
                
                r_data[2859] <= r_data[2858];
                
                r_data[2860] <= r_data[2859];
                
                r_data[2861] <= r_data[2860];
                
                r_data[2862] <= r_data[2861];
                
                r_data[2863] <= r_data[2862];
                
                r_data[2864] <= r_data[2863];
                
                r_data[2865] <= r_data[2864];
                
                r_data[2866] <= r_data[2865];
                
                r_data[2867] <= r_data[2866];
                
                r_data[2868] <= r_data[2867];
                
                r_data[2869] <= r_data[2868];
                
                r_data[2870] <= r_data[2869];
                
                r_data[2871] <= r_data[2870];
                
                r_data[2872] <= r_data[2871];
                
                r_data[2873] <= r_data[2872];
                
                r_data[2874] <= r_data[2873];
                
                r_data[2875] <= r_data[2874];
                
                r_data[2876] <= r_data[2875];
                
                r_data[2877] <= r_data[2876];
                
                r_data[2878] <= r_data[2877];
                
                r_data[2879] <= r_data[2878];
                
                r_data[2880] <= r_data[2879];
                
                r_data[2881] <= r_data[2880];
                
                r_data[2882] <= r_data[2881];
                
                r_data[2883] <= r_data[2882];
                
                r_data[2884] <= r_data[2883];
                
                r_data[2885] <= r_data[2884];
                
                r_data[2886] <= r_data[2885];
                
                r_data[2887] <= r_data[2886];
                
                r_data[2888] <= r_data[2887];
                
                r_data[2889] <= r_data[2888];
                
                r_data[2890] <= r_data[2889];
                
                r_data[2891] <= r_data[2890];
                
                r_data[2892] <= r_data[2891];
                
                r_data[2893] <= r_data[2892];
                
                r_data[2894] <= r_data[2893];
                
                r_data[2895] <= r_data[2894];
                
                r_data[2896] <= r_data[2895];
                
                r_data[2897] <= r_data[2896];
                
                r_data[2898] <= r_data[2897];
                
                r_data[2899] <= r_data[2898];
                
                r_data[2900] <= r_data[2899];
                
                r_data[2901] <= r_data[2900];
                
                r_data[2902] <= r_data[2901];
                
                r_data[2903] <= r_data[2902];
                
                r_data[2904] <= r_data[2903];
                
                r_data[2905] <= r_data[2904];
                
                r_data[2906] <= r_data[2905];
                
                r_data[2907] <= r_data[2906];
                
                r_data[2908] <= r_data[2907];
                
                r_data[2909] <= r_data[2908];
                
                r_data[2910] <= r_data[2909];
                
                r_data[2911] <= r_data[2910];
                
                r_data[2912] <= r_data[2911];
                
                r_data[2913] <= r_data[2912];
                
                r_data[2914] <= r_data[2913];
                
                r_data[2915] <= r_data[2914];
                
                r_data[2916] <= r_data[2915];
                
                r_data[2917] <= r_data[2916];
                
                r_data[2918] <= r_data[2917];
                
                r_data[2919] <= r_data[2918];
                
                r_data[2920] <= r_data[2919];
                
                r_data[2921] <= r_data[2920];
                
                r_data[2922] <= r_data[2921];
                
                r_data[2923] <= r_data[2922];
                
                r_data[2924] <= r_data[2923];
                
                r_data[2925] <= r_data[2924];
                
                r_data[2926] <= r_data[2925];
                
                r_data[2927] <= r_data[2926];
                
                r_data[2928] <= r_data[2927];
                
                r_data[2929] <= r_data[2928];
                
                r_data[2930] <= r_data[2929];
                
                r_data[2931] <= r_data[2930];
                
                r_data[2932] <= r_data[2931];
                
                r_data[2933] <= r_data[2932];
                
                r_data[2934] <= r_data[2933];
                
                r_data[2935] <= r_data[2934];
                
                r_data[2936] <= r_data[2935];
                
                r_data[2937] <= r_data[2936];
                
                r_data[2938] <= r_data[2937];
                
                r_data[2939] <= r_data[2938];
                
                r_data[2940] <= r_data[2939];
                
                r_data[2941] <= r_data[2940];
                
                r_data[2942] <= r_data[2941];
                
                r_data[2943] <= r_data[2942];
                
                r_data[2944] <= r_data[2943];
                
                r_data[2945] <= r_data[2944];
                
                r_data[2946] <= r_data[2945];
                
                r_data[2947] <= r_data[2946];
                
                r_data[2948] <= r_data[2947];
                
                r_data[2949] <= r_data[2948];
                
                r_data[2950] <= r_data[2949];
                
                r_data[2951] <= r_data[2950];
                
                r_data[2952] <= r_data[2951];
                
                r_data[2953] <= r_data[2952];
                
                r_data[2954] <= r_data[2953];
                
                r_data[2955] <= r_data[2954];
                
                r_data[2956] <= r_data[2955];
                
                r_data[2957] <= r_data[2956];
                
                r_data[2958] <= r_data[2957];
                
                r_data[2959] <= r_data[2958];
                
                r_data[2960] <= r_data[2959];
                
                r_data[2961] <= r_data[2960];
                
                r_data[2962] <= r_data[2961];
                
                r_data[2963] <= r_data[2962];
                
                r_data[2964] <= r_data[2963];
                
                r_data[2965] <= r_data[2964];
                
                r_data[2966] <= r_data[2965];
                
                r_data[2967] <= r_data[2966];
                
                r_data[2968] <= r_data[2967];
                
                r_data[2969] <= r_data[2968];
                
                r_data[2970] <= r_data[2969];
                
                r_data[2971] <= r_data[2970];
                
                r_data[2972] <= r_data[2971];
                
                r_data[2973] <= r_data[2972];
                
                r_data[2974] <= r_data[2973];
                
                r_data[2975] <= r_data[2974];
                
                r_data[2976] <= r_data[2975];
                
                r_data[2977] <= r_data[2976];
                
                r_data[2978] <= r_data[2977];
                
                r_data[2979] <= r_data[2978];
                
                r_data[2980] <= r_data[2979];
                
                r_data[2981] <= r_data[2980];
                
                r_data[2982] <= r_data[2981];
                
                r_data[2983] <= r_data[2982];
                
                r_data[2984] <= r_data[2983];
                
                r_data[2985] <= r_data[2984];
                
                r_data[2986] <= r_data[2985];
                
                r_data[2987] <= r_data[2986];
                
                r_data[2988] <= r_data[2987];
                
                r_data[2989] <= r_data[2988];
                
                r_data[2990] <= r_data[2989];
                
                r_data[2991] <= r_data[2990];
                
                r_data[2992] <= r_data[2991];
                
                r_data[2993] <= r_data[2992];
                
                r_data[2994] <= r_data[2993];
                
                r_data[2995] <= r_data[2994];
                
                r_data[2996] <= r_data[2995];
                
                r_data[2997] <= r_data[2996];
                
                r_data[2998] <= r_data[2997];
                
                r_data[2999] <= r_data[2998];
                
                r_data[3000] <= r_data[2999];
                
                r_data[3001] <= r_data[3000];
                
                r_data[3002] <= r_data[3001];
                
                r_data[3003] <= r_data[3002];
                
                r_data[3004] <= r_data[3003];
                
                r_data[3005] <= r_data[3004];
                
                r_data[3006] <= r_data[3005];
                
                r_data[3007] <= r_data[3006];
                
                r_data[3008] <= r_data[3007];
                
                r_data[3009] <= r_data[3008];
                
                r_data[3010] <= r_data[3009];
                
                r_data[3011] <= r_data[3010];
                
                r_data[3012] <= r_data[3011];
                
                r_data[3013] <= r_data[3012];
                
                r_data[3014] <= r_data[3013];
                
                r_data[3015] <= r_data[3014];
                
                r_data[3016] <= r_data[3015];
                
                r_data[3017] <= r_data[3016];
                
                r_data[3018] <= r_data[3017];
                
                r_data[3019] <= r_data[3018];
                
                r_data[3020] <= r_data[3019];
                
                r_data[3021] <= r_data[3020];
                
                r_data[3022] <= r_data[3021];
                
                r_data[3023] <= r_data[3022];
                
                r_data[3024] <= r_data[3023];
                
                r_data[3025] <= r_data[3024];
                
                r_data[3026] <= r_data[3025];
                
                r_data[3027] <= r_data[3026];
                
                r_data[3028] <= r_data[3027];
                
                r_data[3029] <= r_data[3028];
                
                r_data[3030] <= r_data[3029];
                
                r_data[3031] <= r_data[3030];
                
                r_data[3032] <= r_data[3031];
                
                r_data[3033] <= r_data[3032];
                
                r_data[3034] <= r_data[3033];
                
                r_data[3035] <= r_data[3034];
                
                r_data[3036] <= r_data[3035];
                
                r_data[3037] <= r_data[3036];
                
                r_data[3038] <= r_data[3037];
                
                r_data[3039] <= r_data[3038];
                
                r_data[3040] <= r_data[3039];
                
                r_data[3041] <= r_data[3040];
                
                r_data[3042] <= r_data[3041];
                
                r_data[3043] <= r_data[3042];
                
                r_data[3044] <= r_data[3043];
                
                r_data[3045] <= r_data[3044];
                
                r_data[3046] <= r_data[3045];
                
                r_data[3047] <= r_data[3046];
                
                r_data[3048] <= r_data[3047];
                
                r_data[3049] <= r_data[3048];
                
                r_data[3050] <= r_data[3049];
                
                r_data[3051] <= r_data[3050];
                
                r_data[3052] <= r_data[3051];
                
                r_data[3053] <= r_data[3052];
                
                r_data[3054] <= r_data[3053];
                
                r_data[3055] <= r_data[3054];
                
                r_data[3056] <= r_data[3055];
                
                r_data[3057] <= r_data[3056];
                
                r_data[3058] <= r_data[3057];
                
                r_data[3059] <= r_data[3058];
                
                r_data[3060] <= r_data[3059];
                
                r_data[3061] <= r_data[3060];
                
                r_data[3062] <= r_data[3061];
                
                r_data[3063] <= r_data[3062];
                
                r_data[3064] <= r_data[3063];
                
                r_data[3065] <= r_data[3064];
                
                r_data[3066] <= r_data[3065];
                
                r_data[3067] <= r_data[3066];
                
                r_data[3068] <= r_data[3067];
                
                r_data[3069] <= r_data[3068];
                
                r_data[3070] <= r_data[3069];
                
                r_data[3071] <= r_data[3070];
                
                r_data[3072] <= r_data[3071];
                
                r_data[3073] <= r_data[3072];
                
                r_data[3074] <= r_data[3073];
                
                r_data[3075] <= r_data[3074];
                
                r_data[3076] <= r_data[3075];
                
                r_data[3077] <= r_data[3076];
                
                r_data[3078] <= r_data[3077];
                
                r_data[3079] <= r_data[3078];
                
                r_data[3080] <= r_data[3079];
                
                r_data[3081] <= r_data[3080];
                
                r_data[3082] <= r_data[3081];
                
                r_data[3083] <= r_data[3082];
                
                r_data[3084] <= r_data[3083];
                
                r_data[3085] <= r_data[3084];
                
                r_data[3086] <= r_data[3085];
                
                r_data[3087] <= r_data[3086];
                
                r_data[3088] <= r_data[3087];
                
                r_data[3089] <= r_data[3088];
                
                r_data[3090] <= r_data[3089];
                
                r_data[3091] <= r_data[3090];
                
                r_data[3092] <= r_data[3091];
                
                r_data[3093] <= r_data[3092];
                
                r_data[3094] <= r_data[3093];
                
                r_data[3095] <= r_data[3094];
                
                r_data[3096] <= r_data[3095];
                
                r_data[3097] <= r_data[3096];
                
                r_data[3098] <= r_data[3097];
                
                r_data[3099] <= r_data[3098];
                
                r_data[3100] <= r_data[3099];
                
                r_data[3101] <= r_data[3100];
                
                r_data[3102] <= r_data[3101];
                
                r_data[3103] <= r_data[3102];
                
                r_data[3104] <= r_data[3103];
                
                r_data[3105] <= r_data[3104];
                
                r_data[3106] <= r_data[3105];
                
                r_data[3107] <= r_data[3106];
                
                r_data[3108] <= r_data[3107];
                
                r_data[3109] <= r_data[3108];
                
                r_data[3110] <= r_data[3109];
                
                r_data[3111] <= r_data[3110];
                
                r_data[3112] <= r_data[3111];
                
                r_data[3113] <= r_data[3112];
                
                r_data[3114] <= r_data[3113];
                
                r_data[3115] <= r_data[3114];
                
                r_data[3116] <= r_data[3115];
                
                r_data[3117] <= r_data[3116];
                
                r_data[3118] <= r_data[3117];
                
                r_data[3119] <= r_data[3118];
                
                r_data[3120] <= r_data[3119];
                
                r_data[3121] <= r_data[3120];
                
                r_data[3122] <= r_data[3121];
                
                r_data[3123] <= r_data[3122];
                
                r_data[3124] <= r_data[3123];
                
                r_data[3125] <= r_data[3124];
                
                r_data[3126] <= r_data[3125];
                
                r_data[3127] <= r_data[3126];
                
                r_data[3128] <= r_data[3127];
                
                r_data[3129] <= r_data[3128];
                
                r_data[3130] <= r_data[3129];
                
                r_data[3131] <= r_data[3130];
                
                r_data[3132] <= r_data[3131];
                
                r_data[3133] <= r_data[3132];
                
                r_data[3134] <= r_data[3133];
                
                r_data[3135] <= r_data[3134];
                
                r_data[3136] <= r_data[3135];
                
                r_data[3137] <= r_data[3136];
                
                r_data[3138] <= r_data[3137];
                
                r_data[3139] <= r_data[3138];
                
                r_data[3140] <= r_data[3139];
                
                r_data[3141] <= r_data[3140];
                
                r_data[3142] <= r_data[3141];
                
                r_data[3143] <= r_data[3142];
                
                r_data[3144] <= r_data[3143];
                
                r_data[3145] <= r_data[3144];
                
                r_data[3146] <= r_data[3145];
                
                r_data[3147] <= r_data[3146];
                
                r_data[3148] <= r_data[3147];
                
                r_data[3149] <= r_data[3148];
                
                r_data[3150] <= r_data[3149];
                
                r_data[3151] <= r_data[3150];
                
                r_data[3152] <= r_data[3151];
                
                r_data[3153] <= r_data[3152];
                
                r_data[3154] <= r_data[3153];
                
                r_data[3155] <= r_data[3154];
                
                r_data[3156] <= r_data[3155];
                
                r_data[3157] <= r_data[3156];
                
                r_data[3158] <= r_data[3157];
                
                r_data[3159] <= r_data[3158];
                
                r_data[3160] <= r_data[3159];
                
                r_data[3161] <= r_data[3160];
                
                r_data[3162] <= r_data[3161];
                
                r_data[3163] <= r_data[3162];
                
                r_data[3164] <= r_data[3163];
                
                r_data[3165] <= r_data[3164];
                
                r_data[3166] <= r_data[3165];
                
                r_data[3167] <= r_data[3166];
                
                r_data[3168] <= r_data[3167];
                
                r_data[3169] <= r_data[3168];
                
                r_data[3170] <= r_data[3169];
                
                r_data[3171] <= r_data[3170];
                
                r_data[3172] <= r_data[3171];
                
                r_data[3173] <= r_data[3172];
                
                r_data[3174] <= r_data[3173];
                
                r_data[3175] <= r_data[3174];
                
                r_data[3176] <= r_data[3175];
                
                r_data[3177] <= r_data[3176];
                
                r_data[3178] <= r_data[3177];
                
                r_data[3179] <= r_data[3178];
                
                r_data[3180] <= r_data[3179];
                
                r_data[3181] <= r_data[3180];
                
                r_data[3182] <= r_data[3181];
                
                r_data[3183] <= r_data[3182];
                
                r_data[3184] <= r_data[3183];
                
                r_data[3185] <= r_data[3184];
                
                r_data[3186] <= r_data[3185];
                
                r_data[3187] <= r_data[3186];
                
                r_data[3188] <= r_data[3187];
                
                r_data[3189] <= r_data[3188];
                
                r_data[3190] <= r_data[3189];
                
                r_data[3191] <= r_data[3190];
                
                r_data[3192] <= r_data[3191];
                
                r_data[3193] <= r_data[3192];
                
                r_data[3194] <= r_data[3193];
                
                r_data[3195] <= r_data[3194];
                
                r_data[3196] <= r_data[3195];
                
                r_data[3197] <= r_data[3196];
                
                r_data[3198] <= r_data[3197];
                
                r_data[3199] <= r_data[3198];
                
                r_data[3200] <= r_data[3199];
                
                r_data[3201] <= r_data[3200];
                
                r_data[3202] <= r_data[3201];
                
                r_data[3203] <= r_data[3202];
                
                r_data[3204] <= r_data[3203];
                
                r_data[3205] <= r_data[3204];
                
                r_data[3206] <= r_data[3205];
                
                r_data[3207] <= r_data[3206];
                
                r_data[3208] <= r_data[3207];
                
                r_data[3209] <= r_data[3208];
                
                r_data[3210] <= r_data[3209];
                
                r_data[3211] <= r_data[3210];
                
                r_data[3212] <= r_data[3211];
                
                r_data[3213] <= r_data[3212];
                
                r_data[3214] <= r_data[3213];
                
                r_data[3215] <= r_data[3214];
                
                r_data[3216] <= r_data[3215];
                
                r_data[3217] <= r_data[3216];
                
                r_data[3218] <= r_data[3217];
                
                r_data[3219] <= r_data[3218];
                
                r_data[3220] <= r_data[3219];
                
                r_data[3221] <= r_data[3220];
                
                r_data[3222] <= r_data[3221];
                
                r_data[3223] <= r_data[3222];
                
                r_data[3224] <= r_data[3223];
                
                r_data[3225] <= r_data[3224];
                
                r_data[3226] <= r_data[3225];
                
                r_data[3227] <= r_data[3226];
                
                r_data[3228] <= r_data[3227];
                
                r_data[3229] <= r_data[3228];
                
                r_data[3230] <= r_data[3229];
                
                r_data[3231] <= r_data[3230];
                
                r_data[3232] <= r_data[3231];
                
                r_data[3233] <= r_data[3232];
                
                r_data[3234] <= r_data[3233];
                
                r_data[3235] <= r_data[3234];
                
                r_data[3236] <= r_data[3235];
                
                r_data[3237] <= r_data[3236];
                
                r_data[3238] <= r_data[3237];
                
                r_data[3239] <= r_data[3238];
                
                r_data[3240] <= r_data[3239];
                
                r_data[3241] <= r_data[3240];
                
                r_data[3242] <= r_data[3241];
                
                r_data[3243] <= r_data[3242];
                
                r_data[3244] <= r_data[3243];
                
                r_data[3245] <= r_data[3244];
                
                r_data[3246] <= r_data[3245];
                
                r_data[3247] <= r_data[3246];
                
                r_data[3248] <= r_data[3247];
                
                r_data[3249] <= r_data[3248];
                
                r_data[3250] <= r_data[3249];
                
                r_data[3251] <= r_data[3250];
                
                r_data[3252] <= r_data[3251];
                
                r_data[3253] <= r_data[3252];
                
                r_data[3254] <= r_data[3253];
                
                r_data[3255] <= r_data[3254];
                
                r_data[3256] <= r_data[3255];
                
                r_data[3257] <= r_data[3256];
                
                r_data[3258] <= r_data[3257];
                
                r_data[3259] <= r_data[3258];
                
                r_data[3260] <= r_data[3259];
                
                r_data[3261] <= r_data[3260];
                
                r_data[3262] <= r_data[3261];
                
                r_data[3263] <= r_data[3262];
                
                r_data[3264] <= r_data[3263];
                
                r_data[3265] <= r_data[3264];
                
                r_data[3266] <= r_data[3265];
                
                r_data[3267] <= r_data[3266];
                
                r_data[3268] <= r_data[3267];
                
                r_data[3269] <= r_data[3268];
                
                r_data[3270] <= r_data[3269];
                
                r_data[3271] <= r_data[3270];
                
                r_data[3272] <= r_data[3271];
                
                r_data[3273] <= r_data[3272];
                
                r_data[3274] <= r_data[3273];
                
                r_data[3275] <= r_data[3274];
                
                r_data[3276] <= r_data[3275];
                
                r_data[3277] <= r_data[3276];
                
                r_data[3278] <= r_data[3277];
                
                r_data[3279] <= r_data[3278];
                
                r_data[3280] <= r_data[3279];
                
                r_data[3281] <= r_data[3280];
                
                r_data[3282] <= r_data[3281];
                
                r_data[3283] <= r_data[3282];
                
                r_data[3284] <= r_data[3283];
                
                r_data[3285] <= r_data[3284];
                
                r_data[3286] <= r_data[3285];
                
                r_data[3287] <= r_data[3286];
                
                r_data[3288] <= r_data[3287];
                
                r_data[3289] <= r_data[3288];
                
                r_data[3290] <= r_data[3289];
                
                r_data[3291] <= r_data[3290];
                
                r_data[3292] <= r_data[3291];
                
                r_data[3293] <= r_data[3292];
                
                r_data[3294] <= r_data[3293];
                
                r_data[3295] <= r_data[3294];
                
                r_data[3296] <= r_data[3295];
                
                r_data[3297] <= r_data[3296];
                
                r_data[3298] <= r_data[3297];
                
                r_data[3299] <= r_data[3298];
                
                r_data[3300] <= r_data[3299];
                
                r_data[3301] <= r_data[3300];
                
                r_data[3302] <= r_data[3301];
                
                r_data[3303] <= r_data[3302];
                
                r_data[3304] <= r_data[3303];
                
                r_data[3305] <= r_data[3304];
                
                r_data[3306] <= r_data[3305];
                
                r_data[3307] <= r_data[3306];
                
                r_data[3308] <= r_data[3307];
                
                r_data[3309] <= r_data[3308];
                
                r_data[3310] <= r_data[3309];
                
                r_data[3311] <= r_data[3310];
                
                r_data[3312] <= r_data[3311];
                
                r_data[3313] <= r_data[3312];
                
                r_data[3314] <= r_data[3313];
                
                r_data[3315] <= r_data[3314];
                
                r_data[3316] <= r_data[3315];
                
                r_data[3317] <= r_data[3316];
                
                r_data[3318] <= r_data[3317];
                
                r_data[3319] <= r_data[3318];
                
                r_data[3320] <= r_data[3319];
                
                r_data[3321] <= r_data[3320];
                
                r_data[3322] <= r_data[3321];
                
                r_data[3323] <= r_data[3322];
                
                r_data[3324] <= r_data[3323];
                
                r_data[3325] <= r_data[3324];
                
                r_data[3326] <= r_data[3325];
                
                r_data[3327] <= r_data[3326];
                
                r_data[3328] <= r_data[3327];
                
                r_data[3329] <= r_data[3328];
                
                r_data[3330] <= r_data[3329];
                
                r_data[3331] <= r_data[3330];
                
                r_data[3332] <= r_data[3331];
                
                r_data[3333] <= r_data[3332];
                
                r_data[3334] <= r_data[3333];
                
                r_data[3335] <= r_data[3334];
                
                r_data[3336] <= r_data[3335];
                
                r_data[3337] <= r_data[3336];
                
                r_data[3338] <= r_data[3337];
                
                r_data[3339] <= r_data[3338];
                
                r_data[3340] <= r_data[3339];
                
                r_data[3341] <= r_data[3340];
                
                r_data[3342] <= r_data[3341];
                
                r_data[3343] <= r_data[3342];
                
                r_data[3344] <= r_data[3343];
                
                r_data[3345] <= r_data[3344];
                
                r_data[3346] <= r_data[3345];
                
                r_data[3347] <= r_data[3346];
                
                r_data[3348] <= r_data[3347];
                
                r_data[3349] <= r_data[3348];
                
                r_data[3350] <= r_data[3349];
                
                r_data[3351] <= r_data[3350];
                
                r_data[3352] <= r_data[3351];
                
                r_data[3353] <= r_data[3352];
                
                r_data[3354] <= r_data[3353];
                
                r_data[3355] <= r_data[3354];
                
                r_data[3356] <= r_data[3355];
                
                r_data[3357] <= r_data[3356];
                
                r_data[3358] <= r_data[3357];
                
                r_data[3359] <= r_data[3358];
                
                r_data[3360] <= r_data[3359];
                
                r_data[3361] <= r_data[3360];
                
                r_data[3362] <= r_data[3361];
                
                r_data[3363] <= r_data[3362];
                
                r_data[3364] <= r_data[3363];
                
                r_data[3365] <= r_data[3364];
                
                r_data[3366] <= r_data[3365];
                
                r_data[3367] <= r_data[3366];
                
                r_data[3368] <= r_data[3367];
                
                r_data[3369] <= r_data[3368];
                
                r_data[3370] <= r_data[3369];
                
                r_data[3371] <= r_data[3370];
                
                r_data[3372] <= r_data[3371];
                
                r_data[3373] <= r_data[3372];
                
                r_data[3374] <= r_data[3373];
                
                r_data[3375] <= r_data[3374];
                
                r_data[3376] <= r_data[3375];
                
                r_data[3377] <= r_data[3376];
                
                r_data[3378] <= r_data[3377];
                
                r_data[3379] <= r_data[3378];
                
                r_data[3380] <= r_data[3379];
                
                r_data[3381] <= r_data[3380];
                
                r_data[3382] <= r_data[3381];
                
                r_data[3383] <= r_data[3382];
                
                r_data[3384] <= r_data[3383];
                
                r_data[3385] <= r_data[3384];
                
                r_data[3386] <= r_data[3385];
                
                r_data[3387] <= r_data[3386];
                
                r_data[3388] <= r_data[3387];
                
                r_data[3389] <= r_data[3388];
                
                r_data[3390] <= r_data[3389];
                
                r_data[3391] <= r_data[3390];
                
                r_data[3392] <= r_data[3391];
                
                r_data[3393] <= r_data[3392];
                
                r_data[3394] <= r_data[3393];
                
                r_data[3395] <= r_data[3394];
                
                r_data[3396] <= r_data[3395];
                
                r_data[3397] <= r_data[3396];
                
                r_data[3398] <= r_data[3397];
                
                r_data[3399] <= r_data[3398];
                
                r_data[3400] <= r_data[3399];
                
                r_data[3401] <= r_data[3400];
                
                r_data[3402] <= r_data[3401];
                
                r_data[3403] <= r_data[3402];
                
                r_data[3404] <= r_data[3403];
                
                r_data[3405] <= r_data[3404];
                
                r_data[3406] <= r_data[3405];
                
                r_data[3407] <= r_data[3406];
                
                r_data[3408] <= r_data[3407];
                
                r_data[3409] <= r_data[3408];
                
                r_data[3410] <= r_data[3409];
                
                r_data[3411] <= r_data[3410];
                
                r_data[3412] <= r_data[3411];
                
                r_data[3413] <= r_data[3412];
                
                r_data[3414] <= r_data[3413];
                
                r_data[3415] <= r_data[3414];
                
                r_data[3416] <= r_data[3415];
                
                r_data[3417] <= r_data[3416];
                
                r_data[3418] <= r_data[3417];
                
                r_data[3419] <= r_data[3418];
                
                r_data[3420] <= r_data[3419];
                
                r_data[3421] <= r_data[3420];
                
                r_data[3422] <= r_data[3421];
                
                r_data[3423] <= r_data[3422];
                
                r_data[3424] <= r_data[3423];
                
                r_data[3425] <= r_data[3424];
                
                r_data[3426] <= r_data[3425];
                
                r_data[3427] <= r_data[3426];
                
                r_data[3428] <= r_data[3427];
                
                r_data[3429] <= r_data[3428];
                
                r_data[3430] <= r_data[3429];
                
                r_data[3431] <= r_data[3430];
                
                r_data[3432] <= r_data[3431];
                
                r_data[3433] <= r_data[3432];
                
                r_data[3434] <= r_data[3433];
                
                r_data[3435] <= r_data[3434];
                
                r_data[3436] <= r_data[3435];
                
                r_data[3437] <= r_data[3436];
                
                r_data[3438] <= r_data[3437];
                
                r_data[3439] <= r_data[3438];
                
                r_data[3440] <= r_data[3439];
                
                r_data[3441] <= r_data[3440];
                
                r_data[3442] <= r_data[3441];
                
                r_data[3443] <= r_data[3442];
                
                r_data[3444] <= r_data[3443];
                
                r_data[3445] <= r_data[3444];
                
                r_data[3446] <= r_data[3445];
                
                r_data[3447] <= r_data[3446];
                
                r_data[3448] <= r_data[3447];
                
                r_data[3449] <= r_data[3448];
                
                r_data[3450] <= r_data[3449];
                
                r_data[3451] <= r_data[3450];
                
                r_data[3452] <= r_data[3451];
                
                r_data[3453] <= r_data[3452];
                
                r_data[3454] <= r_data[3453];
                
                r_data[3455] <= r_data[3454];
                
                r_data[3456] <= r_data[3455];
                
                r_data[3457] <= r_data[3456];
                
                r_data[3458] <= r_data[3457];
                
                r_data[3459] <= r_data[3458];
                
                r_data[3460] <= r_data[3459];
                
                r_data[3461] <= r_data[3460];
                
                r_data[3462] <= r_data[3461];
                
                r_data[3463] <= r_data[3462];
                
                r_data[3464] <= r_data[3463];
                
                r_data[3465] <= r_data[3464];
                
                r_data[3466] <= r_data[3465];
                
                r_data[3467] <= r_data[3466];
                
                r_data[3468] <= r_data[3467];
                
                r_data[3469] <= r_data[3468];
                
                r_data[3470] <= r_data[3469];
                
                r_data[3471] <= r_data[3470];
                
                r_data[3472] <= r_data[3471];
                
                r_data[3473] <= r_data[3472];
                
                r_data[3474] <= r_data[3473];
                
                r_data[3475] <= r_data[3474];
                
                r_data[3476] <= r_data[3475];
                
                r_data[3477] <= r_data[3476];
                
                r_data[3478] <= r_data[3477];
                
                r_data[3479] <= r_data[3478];
                
                r_data[3480] <= r_data[3479];
                
                r_data[3481] <= r_data[3480];
                
                r_data[3482] <= r_data[3481];
                
                r_data[3483] <= r_data[3482];
                
                r_data[3484] <= r_data[3483];
                
                r_data[3485] <= r_data[3484];
                
                r_data[3486] <= r_data[3485];
                
                r_data[3487] <= r_data[3486];
                
                r_data[3488] <= r_data[3487];
                
                r_data[3489] <= r_data[3488];
                
                r_data[3490] <= r_data[3489];
                
                r_data[3491] <= r_data[3490];
                
                r_data[3492] <= r_data[3491];
                
                r_data[3493] <= r_data[3492];
                
                r_data[3494] <= r_data[3493];
                
                r_data[3495] <= r_data[3494];
                
                r_data[3496] <= r_data[3495];
                
                r_data[3497] <= r_data[3496];
                
                r_data[3498] <= r_data[3497];
                
                r_data[3499] <= r_data[3498];
                
                r_data[3500] <= r_data[3499];
                
                r_data[3501] <= r_data[3500];
                
                r_data[3502] <= r_data[3501];
                
                r_data[3503] <= r_data[3502];
                
                r_data[3504] <= r_data[3503];
                
                r_data[3505] <= r_data[3504];
                
                r_data[3506] <= r_data[3505];
                
                r_data[3507] <= r_data[3506];
                
                r_data[3508] <= r_data[3507];
                
                r_data[3509] <= r_data[3508];
                
                r_data[3510] <= r_data[3509];
                
                r_data[3511] <= r_data[3510];
                
                r_data[3512] <= r_data[3511];
                
                r_data[3513] <= r_data[3512];
                
                r_data[3514] <= r_data[3513];
                
                r_data[3515] <= r_data[3514];
                
                r_data[3516] <= r_data[3515];
                
                r_data[3517] <= r_data[3516];
                
                r_data[3518] <= r_data[3517];
                
                r_data[3519] <= r_data[3518];
                
                r_data[3520] <= r_data[3519];
                
                r_data[3521] <= r_data[3520];
                
                r_data[3522] <= r_data[3521];
                
                r_data[3523] <= r_data[3522];
                
                r_data[3524] <= r_data[3523];
                
                r_data[3525] <= r_data[3524];
                
                r_data[3526] <= r_data[3525];
                
                r_data[3527] <= r_data[3526];
                
                r_data[3528] <= r_data[3527];
                
                r_data[3529] <= r_data[3528];
                
                r_data[3530] <= r_data[3529];
                
                r_data[3531] <= r_data[3530];
                
                r_data[3532] <= r_data[3531];
                
                r_data[3533] <= r_data[3532];
                
                r_data[3534] <= r_data[3533];
                
                r_data[3535] <= r_data[3534];
                
                r_data[3536] <= r_data[3535];
                
                r_data[3537] <= r_data[3536];
                
                r_data[3538] <= r_data[3537];
                
                r_data[3539] <= r_data[3538];
                
                r_data[3540] <= r_data[3539];
                
                r_data[3541] <= r_data[3540];
                
                r_data[3542] <= r_data[3541];
                
                r_data[3543] <= r_data[3542];
                
                r_data[3544] <= r_data[3543];
                
                r_data[3545] <= r_data[3544];
                
                r_data[3546] <= r_data[3545];
                
                r_data[3547] <= r_data[3546];
                
                r_data[3548] <= r_data[3547];
                
                r_data[3549] <= r_data[3548];
                
                r_data[3550] <= r_data[3549];
                
                r_data[3551] <= r_data[3550];
                
                r_data[3552] <= r_data[3551];
                
                r_data[3553] <= r_data[3552];
                
                r_data[3554] <= r_data[3553];
                
                r_data[3555] <= r_data[3554];
                
                r_data[3556] <= r_data[3555];
                
                r_data[3557] <= r_data[3556];
                
                r_data[3558] <= r_data[3557];
                
                r_data[3559] <= r_data[3558];
                
                r_data[3560] <= r_data[3559];
                
                r_data[3561] <= r_data[3560];
                
                r_data[3562] <= r_data[3561];
                
                r_data[3563] <= r_data[3562];
                
                r_data[3564] <= r_data[3563];
                
                r_data[3565] <= r_data[3564];
                
                r_data[3566] <= r_data[3565];
                
                r_data[3567] <= r_data[3566];
                
                r_data[3568] <= r_data[3567];
                
                r_data[3569] <= r_data[3568];
                
                r_data[3570] <= r_data[3569];
                
                r_data[3571] <= r_data[3570];
                
                r_data[3572] <= r_data[3571];
                
                r_data[3573] <= r_data[3572];
                
                r_data[3574] <= r_data[3573];
                
                r_data[3575] <= r_data[3574];
                
                r_data[3576] <= r_data[3575];
                
                r_data[3577] <= r_data[3576];
                
                r_data[3578] <= r_data[3577];
                
                r_data[3579] <= r_data[3578];
                
                r_data[3580] <= r_data[3579];
                
                r_data[3581] <= r_data[3580];
                
                r_data[3582] <= r_data[3581];
                
                r_data[3583] <= r_data[3582];
                
                r_data[3584] <= r_data[3583];
                
                r_data[3585] <= r_data[3584];
                
                r_data[3586] <= r_data[3585];
                
                r_data[3587] <= r_data[3586];
                
                r_data[3588] <= r_data[3587];
                
                r_data[3589] <= r_data[3588];
                
                r_data[3590] <= r_data[3589];
                
                r_data[3591] <= r_data[3590];
                
                r_data[3592] <= r_data[3591];
                
                r_data[3593] <= r_data[3592];
                
                r_data[3594] <= r_data[3593];
                
                r_data[3595] <= r_data[3594];
                
                r_data[3596] <= r_data[3595];
                
                r_data[3597] <= r_data[3596];
                
                r_data[3598] <= r_data[3597];
                
                r_data[3599] <= r_data[3598];
                
                r_data[3600] <= r_data[3599];
                
                r_data[3601] <= r_data[3600];
                
                r_data[3602] <= r_data[3601];
                
                r_data[3603] <= r_data[3602];
                
                r_data[3604] <= r_data[3603];
                
                r_data[3605] <= r_data[3604];
                
                r_data[3606] <= r_data[3605];
                
                r_data[3607] <= r_data[3606];
                
                r_data[3608] <= r_data[3607];
                
                r_data[3609] <= r_data[3608];
                
                r_data[3610] <= r_data[3609];
                
                r_data[3611] <= r_data[3610];
                
                r_data[3612] <= r_data[3611];
                
                r_data[3613] <= r_data[3612];
                
                r_data[3614] <= r_data[3613];
                
                r_data[3615] <= r_data[3614];
                
                r_data[3616] <= r_data[3615];
                
                r_data[3617] <= r_data[3616];
                
                r_data[3618] <= r_data[3617];
                
                r_data[3619] <= r_data[3618];
                
                r_data[3620] <= r_data[3619];
                
                r_data[3621] <= r_data[3620];
                
                r_data[3622] <= r_data[3621];
                
                r_data[3623] <= r_data[3622];
                
                r_data[3624] <= r_data[3623];
                
                r_data[3625] <= r_data[3624];
                
                r_data[3626] <= r_data[3625];
                
                r_data[3627] <= r_data[3626];
                
                r_data[3628] <= r_data[3627];
                
                r_data[3629] <= r_data[3628];
                
                r_data[3630] <= r_data[3629];
                
                r_data[3631] <= r_data[3630];
                
                r_data[3632] <= r_data[3631];
                
                r_data[3633] <= r_data[3632];
                
                r_data[3634] <= r_data[3633];
                
                r_data[3635] <= r_data[3634];
                
                r_data[3636] <= r_data[3635];
                
                r_data[3637] <= r_data[3636];
                
                r_data[3638] <= r_data[3637];
                
                r_data[3639] <= r_data[3638];
                
                r_data[3640] <= r_data[3639];
                
                r_data[3641] <= r_data[3640];
                
                r_data[3642] <= r_data[3641];
                
                r_data[3643] <= r_data[3642];
                
                r_data[3644] <= r_data[3643];
                
                r_data[3645] <= r_data[3644];
                
                r_data[3646] <= r_data[3645];
                
                r_data[3647] <= r_data[3646];
                
                r_data[3648] <= r_data[3647];
                
                r_data[3649] <= r_data[3648];
                
                r_data[3650] <= r_data[3649];
                
                r_data[3651] <= r_data[3650];
                
                r_data[3652] <= r_data[3651];
                
                r_data[3653] <= r_data[3652];
                
                r_data[3654] <= r_data[3653];
                
                r_data[3655] <= r_data[3654];
                
                r_data[3656] <= r_data[3655];
                
                r_data[3657] <= r_data[3656];
                
                r_data[3658] <= r_data[3657];
                
                r_data[3659] <= r_data[3658];
                
                r_data[3660] <= r_data[3659];
                
                r_data[3661] <= r_data[3660];
                
                r_data[3662] <= r_data[3661];
                
                r_data[3663] <= r_data[3662];
                
                r_data[3664] <= r_data[3663];
                
                r_data[3665] <= r_data[3664];
                
                r_data[3666] <= r_data[3665];
                
                r_data[3667] <= r_data[3666];
                
                r_data[3668] <= r_data[3667];
                
                r_data[3669] <= r_data[3668];
                
                r_data[3670] <= r_data[3669];
                
                r_data[3671] <= r_data[3670];
                
                r_data[3672] <= r_data[3671];
                
                r_data[3673] <= r_data[3672];
                
                r_data[3674] <= r_data[3673];
                
                r_data[3675] <= r_data[3674];
                
                r_data[3676] <= r_data[3675];
                
                r_data[3677] <= r_data[3676];
                
                r_data[3678] <= r_data[3677];
                
                r_data[3679] <= r_data[3678];
                
                r_data[3680] <= r_data[3679];
                
                r_data[3681] <= r_data[3680];
                
                r_data[3682] <= r_data[3681];
                
                r_data[3683] <= r_data[3682];
                
                r_data[3684] <= r_data[3683];
                
                r_data[3685] <= r_data[3684];
                
                r_data[3686] <= r_data[3685];
                
                r_data[3687] <= r_data[3686];
                
                r_data[3688] <= r_data[3687];
                
                r_data[3689] <= r_data[3688];
                
                r_data[3690] <= r_data[3689];
                
                r_data[3691] <= r_data[3690];
                
                r_data[3692] <= r_data[3691];
                
                r_data[3693] <= r_data[3692];
                
                r_data[3694] <= r_data[3693];
                
                r_data[3695] <= r_data[3694];
                
                r_data[3696] <= r_data[3695];
                
                r_data[3697] <= r_data[3696];
                
                r_data[3698] <= r_data[3697];
                
                r_data[3699] <= r_data[3698];
                
                r_data[3700] <= r_data[3699];
                
                r_data[3701] <= r_data[3700];
                
                r_data[3702] <= r_data[3701];
                
                r_data[3703] <= r_data[3702];
                
                r_data[3704] <= r_data[3703];
                
                r_data[3705] <= r_data[3704];
                
                r_data[3706] <= r_data[3705];
                
                r_data[3707] <= r_data[3706];
                
                r_data[3708] <= r_data[3707];
                
                r_data[3709] <= r_data[3708];
                
                r_data[3710] <= r_data[3709];
                
                r_data[3711] <= r_data[3710];
                
                r_data[3712] <= r_data[3711];
                
                r_data[3713] <= r_data[3712];
                
                r_data[3714] <= r_data[3713];
                
                r_data[3715] <= r_data[3714];
                
                r_data[3716] <= r_data[3715];
                
                r_data[3717] <= r_data[3716];
                
                r_data[3718] <= r_data[3717];
                
                r_data[3719] <= r_data[3718];
                
                r_data[3720] <= r_data[3719];
                
                r_data[3721] <= r_data[3720];
                
                r_data[3722] <= r_data[3721];
                
                r_data[3723] <= r_data[3722];
                
                r_data[3724] <= r_data[3723];
                
                r_data[3725] <= r_data[3724];
                
                r_data[3726] <= r_data[3725];
                
                r_data[3727] <= r_data[3726];
                
                r_data[3728] <= r_data[3727];
                
                r_data[3729] <= r_data[3728];
                
                r_data[3730] <= r_data[3729];
                
                r_data[3731] <= r_data[3730];
                
                r_data[3732] <= r_data[3731];
                
                r_data[3733] <= r_data[3732];
                
                r_data[3734] <= r_data[3733];
                
                r_data[3735] <= r_data[3734];
                
                r_data[3736] <= r_data[3735];
                
                r_data[3737] <= r_data[3736];
                
                r_data[3738] <= r_data[3737];
                
                r_data[3739] <= r_data[3738];
                
                r_data[3740] <= r_data[3739];
                
                r_data[3741] <= r_data[3740];
                
                r_data[3742] <= r_data[3741];
                
                r_data[3743] <= r_data[3742];
                
                r_data[3744] <= r_data[3743];
                
                r_data[3745] <= r_data[3744];
                
                r_data[3746] <= r_data[3745];
                
                r_data[3747] <= r_data[3746];
                
                r_data[3748] <= r_data[3747];
                
                r_data[3749] <= r_data[3748];
                
                r_data[3750] <= r_data[3749];
                
                r_data[3751] <= r_data[3750];
                
                r_data[3752] <= r_data[3751];
                
                r_data[3753] <= r_data[3752];
                
                r_data[3754] <= r_data[3753];
                
                r_data[3755] <= r_data[3754];
                
                r_data[3756] <= r_data[3755];
                
                r_data[3757] <= r_data[3756];
                
                r_data[3758] <= r_data[3757];
                
                r_data[3759] <= r_data[3758];
                
                r_data[3760] <= r_data[3759];
                
                r_data[3761] <= r_data[3760];
                
                r_data[3762] <= r_data[3761];
                
                r_data[3763] <= r_data[3762];
                
                r_data[3764] <= r_data[3763];
                
                r_data[3765] <= r_data[3764];
                
                r_data[3766] <= r_data[3765];
                
                r_data[3767] <= r_data[3766];
                
                r_data[3768] <= r_data[3767];
                
                r_data[3769] <= r_data[3768];
                
                r_data[3770] <= r_data[3769];
                
                r_data[3771] <= r_data[3770];
                
                r_data[3772] <= r_data[3771];
                
                r_data[3773] <= r_data[3772];
                
                r_data[3774] <= r_data[3773];
                
                r_data[3775] <= r_data[3774];
                
                r_data[3776] <= r_data[3775];
                
                r_data[3777] <= r_data[3776];
                
                r_data[3778] <= r_data[3777];
                
                r_data[3779] <= r_data[3778];
                
                r_data[3780] <= r_data[3779];
                
                r_data[3781] <= r_data[3780];
                
                r_data[3782] <= r_data[3781];
                
                r_data[3783] <= r_data[3782];
                
                r_data[3784] <= r_data[3783];
                
                r_data[3785] <= r_data[3784];
                
                r_data[3786] <= r_data[3785];
                
                r_data[3787] <= r_data[3786];
                
                r_data[3788] <= r_data[3787];
                
                r_data[3789] <= r_data[3788];
                
                r_data[3790] <= r_data[3789];
                
                r_data[3791] <= r_data[3790];
                
                r_data[3792] <= r_data[3791];
                
                r_data[3793] <= r_data[3792];
                
                r_data[3794] <= r_data[3793];
                
                r_data[3795] <= r_data[3794];
                
                r_data[3796] <= r_data[3795];
                
                r_data[3797] <= r_data[3796];
                
                r_data[3798] <= r_data[3797];
                
                r_data[3799] <= r_data[3798];
                
                r_data[3800] <= r_data[3799];
                
                r_data[3801] <= r_data[3800];
                
                r_data[3802] <= r_data[3801];
                
                r_data[3803] <= r_data[3802];
                
                r_data[3804] <= r_data[3803];
                
                r_data[3805] <= r_data[3804];
                
                r_data[3806] <= r_data[3805];
                
                r_data[3807] <= r_data[3806];
                
                r_data[3808] <= r_data[3807];
                
                r_data[3809] <= r_data[3808];
                
                r_data[3810] <= r_data[3809];
                
                r_data[3811] <= r_data[3810];
                
                r_data[3812] <= r_data[3811];
                
                r_data[3813] <= r_data[3812];
                
                r_data[3814] <= r_data[3813];
                
                r_data[3815] <= r_data[3814];
                
                r_data[3816] <= r_data[3815];
                
                r_data[3817] <= r_data[3816];
                
                r_data[3818] <= r_data[3817];
                
                r_data[3819] <= r_data[3818];
                
                r_data[3820] <= r_data[3819];
                
                r_data[3821] <= r_data[3820];
                
                r_data[3822] <= r_data[3821];
                
                r_data[3823] <= r_data[3822];
                
                r_data[3824] <= r_data[3823];
                
                r_data[3825] <= r_data[3824];
                
                r_data[3826] <= r_data[3825];
                
                r_data[3827] <= r_data[3826];
                
                r_data[3828] <= r_data[3827];
                
                r_data[3829] <= r_data[3828];
                
                r_data[3830] <= r_data[3829];
                
                r_data[3831] <= r_data[3830];
                
                r_data[3832] <= r_data[3831];
                
                r_data[3833] <= r_data[3832];
                
                r_data[3834] <= r_data[3833];
                
                r_data[3835] <= r_data[3834];
                
                r_data[3836] <= r_data[3835];
                
                r_data[3837] <= r_data[3836];
                
                r_data[3838] <= r_data[3837];
                
                r_data[3839] <= r_data[3838];
                
                r_data[3840] <= r_data[3839];
                
                r_data[3841] <= r_data[3840];
                
                r_data[3842] <= r_data[3841];
                
                r_data[3843] <= r_data[3842];
                
                r_data[3844] <= r_data[3843];
                
                r_data[3845] <= r_data[3844];
                
                r_data[3846] <= r_data[3845];
                
                r_data[3847] <= r_data[3846];
                
                r_data[3848] <= r_data[3847];
                
                r_data[3849] <= r_data[3848];
                
                r_data[3850] <= r_data[3849];
                
                r_data[3851] <= r_data[3850];
                
                r_data[3852] <= r_data[3851];
                
                r_data[3853] <= r_data[3852];
                
                r_data[3854] <= r_data[3853];
                
                r_data[3855] <= r_data[3854];
                
                r_data[3856] <= r_data[3855];
                
                r_data[3857] <= r_data[3856];
                
                r_data[3858] <= r_data[3857];
                
                r_data[3859] <= r_data[3858];
                
                r_data[3860] <= r_data[3859];
                
                r_data[3861] <= r_data[3860];
                
                r_data[3862] <= r_data[3861];
                
                r_data[3863] <= r_data[3862];
                
                r_data[3864] <= r_data[3863];
                
                r_data[3865] <= r_data[3864];
                
                r_data[3866] <= r_data[3865];
                
                r_data[3867] <= r_data[3866];
                
                r_data[3868] <= r_data[3867];
                
                r_data[3869] <= r_data[3868];
                
                r_data[3870] <= r_data[3869];
                
                r_data[3871] <= r_data[3870];
                
                r_data[3872] <= r_data[3871];
                
                r_data[3873] <= r_data[3872];
                
                r_data[3874] <= r_data[3873];
                
                r_data[3875] <= r_data[3874];
                
                r_data[3876] <= r_data[3875];
                
                r_data[3877] <= r_data[3876];
                
                r_data[3878] <= r_data[3877];
                
                r_data[3879] <= r_data[3878];
                
                r_data[3880] <= r_data[3879];
                
                r_data[3881] <= r_data[3880];
                
                r_data[3882] <= r_data[3881];
                
                r_data[3883] <= r_data[3882];
                
                r_data[3884] <= r_data[3883];
                
                r_data[3885] <= r_data[3884];
                
                r_data[3886] <= r_data[3885];
                
                r_data[3887] <= r_data[3886];
                
                r_data[3888] <= r_data[3887];
                
                r_data[3889] <= r_data[3888];
                
                r_data[3890] <= r_data[3889];
                
                r_data[3891] <= r_data[3890];
                
                r_data[3892] <= r_data[3891];
                
                r_data[3893] <= r_data[3892];
                
                r_data[3894] <= r_data[3893];
                
                r_data[3895] <= r_data[3894];
                
                r_data[3896] <= r_data[3895];
                
                r_data[3897] <= r_data[3896];
                
                r_data[3898] <= r_data[3897];
                
                r_data[3899] <= r_data[3898];
                
                r_data[3900] <= r_data[3899];
                
                r_data[3901] <= r_data[3900];
                
                r_data[3902] <= r_data[3901];
                
                r_data[3903] <= r_data[3902];
                
                r_data[3904] <= r_data[3903];
                
                r_data[3905] <= r_data[3904];
                
                r_data[3906] <= r_data[3905];
                
                r_data[3907] <= r_data[3906];
                
                r_data[3908] <= r_data[3907];
                
                r_data[3909] <= r_data[3908];
                
                r_data[3910] <= r_data[3909];
                
                r_data[3911] <= r_data[3910];
                
                r_data[3912] <= r_data[3911];
                
                r_data[3913] <= r_data[3912];
                
                r_data[3914] <= r_data[3913];
                
                r_data[3915] <= r_data[3914];
                
                r_data[3916] <= r_data[3915];
                
                r_data[3917] <= r_data[3916];
                
                r_data[3918] <= r_data[3917];
                
                r_data[3919] <= r_data[3918];
                
                r_data[3920] <= r_data[3919];
                
                r_data[3921] <= r_data[3920];
                
                r_data[3922] <= r_data[3921];
                
                r_data[3923] <= r_data[3922];
                
                r_data[3924] <= r_data[3923];
                
                r_data[3925] <= r_data[3924];
                
                r_data[3926] <= r_data[3925];
                
                r_data[3927] <= r_data[3926];
                
                r_data[3928] <= r_data[3927];
                
                r_data[3929] <= r_data[3928];
                
                r_data[3930] <= r_data[3929];
                
                r_data[3931] <= r_data[3930];
                
                r_data[3932] <= r_data[3931];
                
                r_data[3933] <= r_data[3932];
                
                r_data[3934] <= r_data[3933];
                
                r_data[3935] <= r_data[3934];
                
                r_data[3936] <= r_data[3935];
                
                r_data[3937] <= r_data[3936];
                
                r_data[3938] <= r_data[3937];
                
                r_data[3939] <= r_data[3938];
                
                r_data[3940] <= r_data[3939];
                
                r_data[3941] <= r_data[3940];
                
                r_data[3942] <= r_data[3941];
                
                r_data[3943] <= r_data[3942];
                
                r_data[3944] <= r_data[3943];
                
                r_data[3945] <= r_data[3944];
                
                r_data[3946] <= r_data[3945];
                
                r_data[3947] <= r_data[3946];
                
                r_data[3948] <= r_data[3947];
                
                r_data[3949] <= r_data[3948];
                
                r_data[3950] <= r_data[3949];
                
                r_data[3951] <= r_data[3950];
                
                r_data[3952] <= r_data[3951];
                
                r_data[3953] <= r_data[3952];
                
                r_data[3954] <= r_data[3953];
                
                r_data[3955] <= r_data[3954];
                
                r_data[3956] <= r_data[3955];
                
                r_data[3957] <= r_data[3956];
                
                r_data[3958] <= r_data[3957];
                
                r_data[3959] <= r_data[3958];
                
                r_data[3960] <= r_data[3959];
                
                r_data[3961] <= r_data[3960];
                
                r_data[3962] <= r_data[3961];
                
                r_data[3963] <= r_data[3962];
                
                r_data[3964] <= r_data[3963];
                
                r_data[3965] <= r_data[3964];
                
                r_data[3966] <= r_data[3965];
                
                r_data[3967] <= r_data[3966];
                
                r_data[3968] <= r_data[3967];
                
                r_data[3969] <= r_data[3968];
                
                r_data[3970] <= r_data[3969];
                
                r_data[3971] <= r_data[3970];
                
                r_data[3972] <= r_data[3971];
                
                r_data[3973] <= r_data[3972];
                
                r_data[3974] <= r_data[3973];
                
                r_data[3975] <= r_data[3974];
                
                r_data[3976] <= r_data[3975];
                
                r_data[3977] <= r_data[3976];
                
                r_data[3978] <= r_data[3977];
                
                r_data[3979] <= r_data[3978];
                
                r_data[3980] <= r_data[3979];
                
                r_data[3981] <= r_data[3980];
                
                r_data[3982] <= r_data[3981];
                
                r_data[3983] <= r_data[3982];
                
                r_data[3984] <= r_data[3983];
                
                r_data[3985] <= r_data[3984];
                
                r_data[3986] <= r_data[3985];
                
                r_data[3987] <= r_data[3986];
                
                r_data[3988] <= r_data[3987];
                
                r_data[3989] <= r_data[3988];
                
                r_data[3990] <= r_data[3989];
                
                r_data[3991] <= r_data[3990];
                
                r_data[3992] <= r_data[3991];
                
                r_data[3993] <= r_data[3992];
                
                r_data[3994] <= r_data[3993];
                
                r_data[3995] <= r_data[3994];
                
                r_data[3996] <= r_data[3995];
                
                r_data[3997] <= r_data[3996];
                
                r_data[3998] <= r_data[3997];
                
                r_data[3999] <= r_data[3998];
                
                r_data[4000] <= r_data[3999];
                
                r_data[4001] <= r_data[4000];
                
                r_data[4002] <= r_data[4001];
                
                r_data[4003] <= r_data[4002];
                
                r_data[4004] <= r_data[4003];
                
                r_data[4005] <= r_data[4004];
                
                r_data[4006] <= r_data[4005];
                
                r_data[4007] <= r_data[4006];
                
                r_data[4008] <= r_data[4007];
                
                r_data[4009] <= r_data[4008];
                
                r_data[4010] <= r_data[4009];
                
                r_data[4011] <= r_data[4010];
                
                r_data[4012] <= r_data[4011];
                
                r_data[4013] <= r_data[4012];
                
                r_data[4014] <= r_data[4013];
                
                r_data[4015] <= r_data[4014];
                
                r_data[4016] <= r_data[4015];
                
                r_data[4017] <= r_data[4016];
                
                r_data[4018] <= r_data[4017];
                
                r_data[4019] <= r_data[4018];
                
                r_data[4020] <= r_data[4019];
                
                r_data[4021] <= r_data[4020];
                
                r_data[4022] <= r_data[4021];
                
                r_data[4023] <= r_data[4022];
                
                r_data[4024] <= r_data[4023];
                
                r_data[4025] <= r_data[4024];
                
                r_data[4026] <= r_data[4025];
                
                r_data[4027] <= r_data[4026];
                
                r_data[4028] <= r_data[4027];
                
                r_data[4029] <= r_data[4028];
                
                r_data[4030] <= r_data[4029];
                
                r_data[4031] <= r_data[4030];
                
                r_data[4032] <= r_data[4031];
                
                r_data[4033] <= r_data[4032];
                
                r_data[4034] <= r_data[4033];
                
                r_data[4035] <= r_data[4034];
                
                r_data[4036] <= r_data[4035];
                
                r_data[4037] <= r_data[4036];
                
                r_data[4038] <= r_data[4037];
                
                r_data[4039] <= r_data[4038];
                
                r_data[4040] <= r_data[4039];
                
                r_data[4041] <= r_data[4040];
                
                r_data[4042] <= r_data[4041];
                
                r_data[4043] <= r_data[4042];
                
                r_data[4044] <= r_data[4043];
                
                r_data[4045] <= r_data[4044];
                
                r_data[4046] <= r_data[4045];
                
                r_data[4047] <= r_data[4046];
                
                r_data[4048] <= r_data[4047];
                
                r_data[4049] <= r_data[4048];
                
                r_data[4050] <= r_data[4049];
                
                r_data[4051] <= r_data[4050];
                
                r_data[4052] <= r_data[4051];
                
                r_data[4053] <= r_data[4052];
                
                r_data[4054] <= r_data[4053];
                
                r_data[4055] <= r_data[4054];
                
                r_data[4056] <= r_data[4055];
                
                r_data[4057] <= r_data[4056];
                
                r_data[4058] <= r_data[4057];
                
                r_data[4059] <= r_data[4058];
                
                r_data[4060] <= r_data[4059];
                
                r_data[4061] <= r_data[4060];
                
                r_data[4062] <= r_data[4061];
                
                r_data[4063] <= r_data[4062];
                
                r_data[4064] <= r_data[4063];
                
                r_data[4065] <= r_data[4064];
                
                r_data[4066] <= r_data[4065];
                
                r_data[4067] <= r_data[4066];
                
                r_data[4068] <= r_data[4067];
                
                r_data[4069] <= r_data[4068];
                
                r_data[4070] <= r_data[4069];
                
                r_data[4071] <= r_data[4070];
                
                r_data[4072] <= r_data[4071];
                
                r_data[4073] <= r_data[4072];
                
                r_data[4074] <= r_data[4073];
                
                r_data[4075] <= r_data[4074];
                
                r_data[4076] <= r_data[4075];
                
                r_data[4077] <= r_data[4076];
                
                r_data[4078] <= r_data[4077];
                
                r_data[4079] <= r_data[4078];
                
                r_data[4080] <= r_data[4079];
                
                r_data[4081] <= r_data[4080];
                
                r_data[4082] <= r_data[4081];
                
                r_data[4083] <= r_data[4082];
                
                r_data[4084] <= r_data[4083];
                
                r_data[4085] <= r_data[4084];
                
                r_data[4086] <= r_data[4085];
                
                r_data[4087] <= r_data[4086];
                
                r_data[4088] <= r_data[4087];
                
                r_data[4089] <= r_data[4088];
                
                r_data[4090] <= r_data[4089];
                
                r_data[4091] <= r_data[4090];
                
                r_data[4092] <= r_data[4091];
                
                r_data[4093] <= r_data[4092];
                
                r_data[4094] <= r_data[4093];
                
                r_data[4095] <= r_data[4094];
                
                r_data[4096] <= r_data[4095];
                
                r_data[4097] <= r_data[4096];
                
                r_data[4098] <= r_data[4097];
                
                r_data[4099] <= r_data[4098];
                
                r_data[4100] <= r_data[4099];
                
                r_data[4101] <= r_data[4100];
                
                r_data[4102] <= r_data[4101];
                
                r_data[4103] <= r_data[4102];
                
                r_data[4104] <= r_data[4103];
                
                r_data[4105] <= r_data[4104];
                
                r_data[4106] <= r_data[4105];
                
                r_data[4107] <= r_data[4106];
                
                r_data[4108] <= r_data[4107];
                
                r_data[4109] <= r_data[4108];
                
                r_data[4110] <= r_data[4109];
                
                r_data[4111] <= r_data[4110];
                
                r_data[4112] <= r_data[4111];
                
                r_data[4113] <= r_data[4112];
                
                r_data[4114] <= r_data[4113];
                
                r_data[4115] <= r_data[4114];
                
                r_data[4116] <= r_data[4115];
                
                r_data[4117] <= r_data[4116];
                
                r_data[4118] <= r_data[4117];
                
                r_data[4119] <= r_data[4118];
                
                r_data[4120] <= r_data[4119];
                
                r_data[4121] <= r_data[4120];
                
                r_data[4122] <= r_data[4121];
                
                r_data[4123] <= r_data[4122];
                
                r_data[4124] <= r_data[4123];
                
                r_data[4125] <= r_data[4124];
                
                r_data[4126] <= r_data[4125];
                
                r_data[4127] <= r_data[4126];
                
                r_data[4128] <= r_data[4127];
                
                r_data[4129] <= r_data[4128];
                
                r_data[4130] <= r_data[4129];
                
                r_data[4131] <= r_data[4130];
                
                r_data[4132] <= r_data[4131];
                
                r_data[4133] <= r_data[4132];
                
                r_data[4134] <= r_data[4133];
                
                r_data[4135] <= r_data[4134];
                
                r_data[4136] <= r_data[4135];
                
                r_data[4137] <= r_data[4136];
                
                r_data[4138] <= r_data[4137];
                
                r_data[4139] <= r_data[4138];
                
                r_data[4140] <= r_data[4139];
                
                r_data[4141] <= r_data[4140];
                
                r_data[4142] <= r_data[4141];
                
                r_data[4143] <= r_data[4142];
                
                r_data[4144] <= r_data[4143];
                
                r_data[4145] <= r_data[4144];
                
                r_data[4146] <= r_data[4145];
                
                r_data[4147] <= r_data[4146];
                
                r_data[4148] <= r_data[4147];
                
                r_data[4149] <= r_data[4148];
                
                r_data[4150] <= r_data[4149];
                
                r_data[4151] <= r_data[4150];
                
                r_data[4152] <= r_data[4151];
                
                r_data[4153] <= r_data[4152];
                
                r_data[4154] <= r_data[4153];
                
                r_data[4155] <= r_data[4154];
                
                r_data[4156] <= r_data[4155];
                
                r_data[4157] <= r_data[4156];
                
                r_data[4158] <= r_data[4157];
                
                r_data[4159] <= r_data[4158];
                
                r_data[4160] <= r_data[4159];
                
                r_data[4161] <= r_data[4160];
                
                r_data[4162] <= r_data[4161];
                
                r_data[4163] <= r_data[4162];
                
                r_data[4164] <= r_data[4163];
                
                r_data[4165] <= r_data[4164];
                
                r_data[4166] <= r_data[4165];
                
                r_data[4167] <= r_data[4166];
                
                r_data[4168] <= r_data[4167];
                
                r_data[4169] <= r_data[4168];
                
                r_data[4170] <= r_data[4169];
                
                r_data[4171] <= r_data[4170];
                
                r_data[4172] <= r_data[4171];
                
                r_data[4173] <= r_data[4172];
                
                r_data[4174] <= r_data[4173];
                
                r_data[4175] <= r_data[4174];
                
                r_data[4176] <= r_data[4175];
                
                r_data[4177] <= r_data[4176];
                
                r_data[4178] <= r_data[4177];
                
                r_data[4179] <= r_data[4178];
                
                r_data[4180] <= r_data[4179];
                
                r_data[4181] <= r_data[4180];
                
                r_data[4182] <= r_data[4181];
                
                r_data[4183] <= r_data[4182];
                
                r_data[4184] <= r_data[4183];
                
                r_data[4185] <= r_data[4184];
                
                r_data[4186] <= r_data[4185];
                
                r_data[4187] <= r_data[4186];
                
                r_data[4188] <= r_data[4187];
                
                r_data[4189] <= r_data[4188];
                
                r_data[4190] <= r_data[4189];
                
                r_data[4191] <= r_data[4190];
                
                r_data[4192] <= r_data[4191];
                
                r_data[4193] <= r_data[4192];
                
                r_data[4194] <= r_data[4193];
                
                r_data[4195] <= r_data[4194];
                
                r_data[4196] <= r_data[4195];
                
                r_data[4197] <= r_data[4196];
                
                r_data[4198] <= r_data[4197];
                
                r_data[4199] <= r_data[4198];
                
                r_data[4200] <= r_data[4199];
                
                r_data[4201] <= r_data[4200];
                
                r_data[4202] <= r_data[4201];
                
                r_data[4203] <= r_data[4202];
                
                r_data[4204] <= r_data[4203];
                
                r_data[4205] <= r_data[4204];
                
                r_data[4206] <= r_data[4205];
                
                r_data[4207] <= r_data[4206];
                
                r_data[4208] <= r_data[4207];
                
                r_data[4209] <= r_data[4208];
                
                r_data[4210] <= r_data[4209];
                
                r_data[4211] <= r_data[4210];
                
                r_data[4212] <= r_data[4211];
                
                r_data[4213] <= r_data[4212];
                
                r_data[4214] <= r_data[4213];
                
                r_data[4215] <= r_data[4214];
                
                r_data[4216] <= r_data[4215];
                
                r_data[4217] <= r_data[4216];
                
                r_data[4218] <= r_data[4217];
                
                r_data[4219] <= r_data[4218];
                
                r_data[4220] <= r_data[4219];
                
                r_data[4221] <= r_data[4220];
                
                r_data[4222] <= r_data[4221];
                
                r_data[4223] <= r_data[4222];
                
                r_data[4224] <= r_data[4223];
                
                r_data[4225] <= r_data[4224];
                
                r_data[4226] <= r_data[4225];
                
                r_data[4227] <= r_data[4226];
                
                r_data[4228] <= r_data[4227];
                
                r_data[4229] <= r_data[4228];
                
                r_data[4230] <= r_data[4229];
                
                r_data[4231] <= r_data[4230];
                
                r_data[4232] <= r_data[4231];
                
                r_data[4233] <= r_data[4232];
                
                r_data[4234] <= r_data[4233];
                
                r_data[4235] <= r_data[4234];
                
                r_data[4236] <= r_data[4235];
                
                r_data[4237] <= r_data[4236];
                
                r_data[4238] <= r_data[4237];
                
                r_data[4239] <= r_data[4238];
                
                r_data[4240] <= r_data[4239];
                
                r_data[4241] <= r_data[4240];
                
                r_data[4242] <= r_data[4241];
                
                r_data[4243] <= r_data[4242];
                
                r_data[4244] <= r_data[4243];
                
                r_data[4245] <= r_data[4244];
                
                r_data[4246] <= r_data[4245];
                
                r_data[4247] <= r_data[4246];
                
                r_data[4248] <= r_data[4247];
                
                r_data[4249] <= r_data[4248];
                
                r_data[4250] <= r_data[4249];
                
                r_data[4251] <= r_data[4250];
                
                r_data[4252] <= r_data[4251];
                
                r_data[4253] <= r_data[4252];
                
                r_data[4254] <= r_data[4253];
                
                r_data[4255] <= r_data[4254];
                
                r_data[4256] <= r_data[4255];
                
                r_data[4257] <= r_data[4256];
                
                r_data[4258] <= r_data[4257];
                
                r_data[4259] <= r_data[4258];
                
                r_data[4260] <= r_data[4259];
                
                r_data[4261] <= r_data[4260];
                
                r_data[4262] <= r_data[4261];
                
                r_data[4263] <= r_data[4262];
                
                r_data[4264] <= r_data[4263];
                
                r_data[4265] <= r_data[4264];
                
                r_data[4266] <= r_data[4265];
                
                r_data[4267] <= r_data[4266];
                
                r_data[4268] <= r_data[4267];
                
                r_data[4269] <= r_data[4268];
                
                r_data[4270] <= r_data[4269];
                
                r_data[4271] <= r_data[4270];
                
                r_data[4272] <= r_data[4271];
                
                r_data[4273] <= r_data[4272];
                
                r_data[4274] <= r_data[4273];
                
                r_data[4275] <= r_data[4274];
                
                r_data[4276] <= r_data[4275];
                
                r_data[4277] <= r_data[4276];
                
                r_data[4278] <= r_data[4277];
                
                r_data[4279] <= r_data[4278];
                
                r_data[4280] <= r_data[4279];
                
                r_data[4281] <= r_data[4280];
                
                r_data[4282] <= r_data[4281];
                
                r_data[4283] <= r_data[4282];
                
                r_data[4284] <= r_data[4283];
                
                r_data[4285] <= r_data[4284];
                
                r_data[4286] <= r_data[4285];
                
                r_data[4287] <= r_data[4286];
                
                r_data[4288] <= r_data[4287];
                
                r_data[4289] <= r_data[4288];
                
                r_data[4290] <= r_data[4289];
                
                r_data[4291] <= r_data[4290];
                
                r_data[4292] <= r_data[4291];
                
                r_data[4293] <= r_data[4292];
                
                r_data[4294] <= r_data[4293];
                
                r_data[4295] <= r_data[4294];
                
                r_data[4296] <= r_data[4295];
                
                r_data[4297] <= r_data[4296];
                
                r_data[4298] <= r_data[4297];
                
                r_data[4299] <= r_data[4298];
                
                r_data[4300] <= r_data[4299];
                
                r_data[4301] <= r_data[4300];
                
                r_data[4302] <= r_data[4301];
                
                r_data[4303] <= r_data[4302];
                
                r_data[4304] <= r_data[4303];
                
                r_data[4305] <= r_data[4304];
                
                r_data[4306] <= r_data[4305];
                
                r_data[4307] <= r_data[4306];
                
                r_data[4308] <= r_data[4307];
                
                r_data[4309] <= r_data[4308];
                
                r_data[4310] <= r_data[4309];
                
                r_data[4311] <= r_data[4310];
                
                r_data[4312] <= r_data[4311];
                
                r_data[4313] <= r_data[4312];
                
                r_data[4314] <= r_data[4313];
                
                r_data[4315] <= r_data[4314];
                
                r_data[4316] <= r_data[4315];
                
                r_data[4317] <= r_data[4316];
                
                r_data[4318] <= r_data[4317];
                
                r_data[4319] <= r_data[4318];
                
                r_data[4320] <= r_data[4319];
                
                r_data[4321] <= r_data[4320];
                
                r_data[4322] <= r_data[4321];
                
                r_data[4323] <= r_data[4322];
                
                r_data[4324] <= r_data[4323];
                
                r_data[4325] <= r_data[4324];
                
                r_data[4326] <= r_data[4325];
                
                r_data[4327] <= r_data[4326];
                
                r_data[4328] <= r_data[4327];
                
                r_data[4329] <= r_data[4328];
                
                r_data[4330] <= r_data[4329];
                
                r_data[4331] <= r_data[4330];
                
                r_data[4332] <= r_data[4331];
                
                r_data[4333] <= r_data[4332];
                
                r_data[4334] <= r_data[4333];
                
                r_data[4335] <= r_data[4334];
                
                r_data[4336] <= r_data[4335];
                
                r_data[4337] <= r_data[4336];
                
                r_data[4338] <= r_data[4337];
                
                r_data[4339] <= r_data[4338];
                
                r_data[4340] <= r_data[4339];
                
                r_data[4341] <= r_data[4340];
                
                r_data[4342] <= r_data[4341];
                
                r_data[4343] <= r_data[4342];
                
                r_data[4344] <= r_data[4343];
                
                r_data[4345] <= r_data[4344];
                
                r_data[4346] <= r_data[4345];
                
                r_data[4347] <= r_data[4346];
                
                r_data[4348] <= r_data[4347];
                
                r_data[4349] <= r_data[4348];
                
                r_data[4350] <= r_data[4349];
                
                r_data[4351] <= r_data[4350];
                
                r_data[4352] <= r_data[4351];
                
                r_data[4353] <= r_data[4352];
                
                r_data[4354] <= r_data[4353];
                
                r_data[4355] <= r_data[4354];
                
                r_data[4356] <= r_data[4355];
                
                r_data[4357] <= r_data[4356];
                
                r_data[4358] <= r_data[4357];
                
                r_data[4359] <= r_data[4358];
                
                r_data[4360] <= r_data[4359];
                
                r_data[4361] <= r_data[4360];
                
                r_data[4362] <= r_data[4361];
                
                r_data[4363] <= r_data[4362];
                
                r_data[4364] <= r_data[4363];
                
                r_data[4365] <= r_data[4364];
                
                r_data[4366] <= r_data[4365];
                
                r_data[4367] <= r_data[4366];
                
                r_data[4368] <= r_data[4367];
                
                r_data[4369] <= r_data[4368];
                
                r_data[4370] <= r_data[4369];
                
                r_data[4371] <= r_data[4370];
                
                r_data[4372] <= r_data[4371];
                
                r_data[4373] <= r_data[4372];
                
                r_data[4374] <= r_data[4373];
                
                r_data[4375] <= r_data[4374];
                
                r_data[4376] <= r_data[4375];
                
                r_data[4377] <= r_data[4376];
                
                r_data[4378] <= r_data[4377];
                
                r_data[4379] <= r_data[4378];
                
                r_data[4380] <= r_data[4379];
                
                r_data[4381] <= r_data[4380];
                
                r_data[4382] <= r_data[4381];
                
                r_data[4383] <= r_data[4382];
                
                r_data[4384] <= r_data[4383];
                
                r_data[4385] <= r_data[4384];
                
                r_data[4386] <= r_data[4385];
                
                r_data[4387] <= r_data[4386];
                
                r_data[4388] <= r_data[4387];
                
                r_data[4389] <= r_data[4388];
                
                r_data[4390] <= r_data[4389];
                
                r_data[4391] <= r_data[4390];
                
                r_data[4392] <= r_data[4391];
                
                r_data[4393] <= r_data[4392];
                
                r_data[4394] <= r_data[4393];
                
                r_data[4395] <= r_data[4394];
                
                r_data[4396] <= r_data[4395];
                
                r_data[4397] <= r_data[4396];
                
                r_data[4398] <= r_data[4397];
                
                r_data[4399] <= r_data[4398];
                
                r_data[4400] <= r_data[4399];
                
                r_data[4401] <= r_data[4400];
                
                r_data[4402] <= r_data[4401];
                
                r_data[4403] <= r_data[4402];
                
                r_data[4404] <= r_data[4403];
                
                r_data[4405] <= r_data[4404];
                
                r_data[4406] <= r_data[4405];
                
                r_data[4407] <= r_data[4406];
                
                r_data[4408] <= r_data[4407];
                
                r_data[4409] <= r_data[4408];
                
                r_data[4410] <= r_data[4409];
                
                r_data[4411] <= r_data[4410];
                
                r_data[4412] <= r_data[4411];
                
                r_data[4413] <= r_data[4412];
                
                r_data[4414] <= r_data[4413];
                
                r_data[4415] <= r_data[4414];
                
                r_data[4416] <= r_data[4415];
                
                r_data[4417] <= r_data[4416];
                
                r_data[4418] <= r_data[4417];
                
                r_data[4419] <= r_data[4418];
                
                r_data[4420] <= r_data[4419];
                
                r_data[4421] <= r_data[4420];
                
                r_data[4422] <= r_data[4421];
                
                r_data[4423] <= r_data[4422];
                
                r_data[4424] <= r_data[4423];
                
                r_data[4425] <= r_data[4424];
                
                r_data[4426] <= r_data[4425];
                
                r_data[4427] <= r_data[4426];
                
                r_data[4428] <= r_data[4427];
                
                r_data[4429] <= r_data[4428];
                
                r_data[4430] <= r_data[4429];
                
                r_data[4431] <= r_data[4430];
                
                r_data[4432] <= r_data[4431];
                
                r_data[4433] <= r_data[4432];
                
                r_data[4434] <= r_data[4433];
                
                r_data[4435] <= r_data[4434];
                
                r_data[4436] <= r_data[4435];
                
                r_data[4437] <= r_data[4436];
                
                r_data[4438] <= r_data[4437];
                
                r_data[4439] <= r_data[4438];
                
                r_data[4440] <= r_data[4439];
                
                r_data[4441] <= r_data[4440];
                
                r_data[4442] <= r_data[4441];
                
                r_data[4443] <= r_data[4442];
                
                r_data[4444] <= r_data[4443];
                
                r_data[4445] <= r_data[4444];
                
                r_data[4446] <= r_data[4445];
                
                r_data[4447] <= r_data[4446];
                
                r_data[4448] <= r_data[4447];
                
                r_data[4449] <= r_data[4448];
                
                r_data[4450] <= r_data[4449];
                
                r_data[4451] <= r_data[4450];
                
                r_data[4452] <= r_data[4451];
                
                r_data[4453] <= r_data[4452];
                
                r_data[4454] <= r_data[4453];
                
                r_data[4455] <= r_data[4454];
                
                r_data[4456] <= r_data[4455];
                
                r_data[4457] <= r_data[4456];
                
                r_data[4458] <= r_data[4457];
                
                r_data[4459] <= r_data[4458];
                
                r_data[4460] <= r_data[4459];
                
                r_data[4461] <= r_data[4460];
                
                r_data[4462] <= r_data[4461];
                
                r_data[4463] <= r_data[4462];
                
                r_data[4464] <= r_data[4463];
                
                r_data[4465] <= r_data[4464];
                
                r_data[4466] <= r_data[4465];
                
                r_data[4467] <= r_data[4466];
                
                r_data[4468] <= r_data[4467];
                
                r_data[4469] <= r_data[4468];
                
                r_data[4470] <= r_data[4469];
                
                r_data[4471] <= r_data[4470];
                
                r_data[4472] <= r_data[4471];
                
                r_data[4473] <= r_data[4472];
                
                r_data[4474] <= r_data[4473];
                
                r_data[4475] <= r_data[4474];
                
                r_data[4476] <= r_data[4475];
                
                r_data[4477] <= r_data[4476];
                
                r_data[4478] <= r_data[4477];
                
                r_data[4479] <= r_data[4478];
                
                r_data[4480] <= r_data[4479];
                
                r_data[4481] <= r_data[4480];
                
                r_data[4482] <= r_data[4481];
                
                r_data[4483] <= r_data[4482];
                
                r_data[4484] <= r_data[4483];
                
                r_data[4485] <= r_data[4484];
                
                r_data[4486] <= r_data[4485];
                
                r_data[4487] <= r_data[4486];
                
                r_data[4488] <= r_data[4487];
                
                r_data[4489] <= r_data[4488];
                
                r_data[4490] <= r_data[4489];
                
                r_data[4491] <= r_data[4490];
                
                r_data[4492] <= r_data[4491];
                
                r_data[4493] <= r_data[4492];
                
                r_data[4494] <= r_data[4493];
                
                r_data[4495] <= r_data[4494];
                
                r_data[4496] <= r_data[4495];
                
                r_data[4497] <= r_data[4496];
                
                r_data[4498] <= r_data[4497];
                
                r_data[4499] <= r_data[4498];
                
                r_data[4500] <= r_data[4499];
                
                r_data[4501] <= r_data[4500];
                
                r_data[4502] <= r_data[4501];
                
                r_data[4503] <= r_data[4502];
                
                r_data[4504] <= r_data[4503];
                
                r_data[4505] <= r_data[4504];
                
                r_data[4506] <= r_data[4505];
                
                r_data[4507] <= r_data[4506];
                
                r_data[4508] <= r_data[4507];
                
                r_data[4509] <= r_data[4508];
                
                r_data[4510] <= r_data[4509];
                
                r_data[4511] <= r_data[4510];
                
                r_data[4512] <= r_data[4511];
                
                r_data[4513] <= r_data[4512];
                
                r_data[4514] <= r_data[4513];
                
                r_data[4515] <= r_data[4514];
                
                r_data[4516] <= r_data[4515];
                
                r_data[4517] <= r_data[4516];
                
                r_data[4518] <= r_data[4517];
                
                r_data[4519] <= r_data[4518];
                
                r_data[4520] <= r_data[4519];
                
                r_data[4521] <= r_data[4520];
                
                r_data[4522] <= r_data[4521];
                
                r_data[4523] <= r_data[4522];
                
                r_data[4524] <= r_data[4523];
                
                r_data[4525] <= r_data[4524];
                
                r_data[4526] <= r_data[4525];
                
                r_data[4527] <= r_data[4526];
                
                r_data[4528] <= r_data[4527];
                
                r_data[4529] <= r_data[4528];
                
                r_data[4530] <= r_data[4529];
                
                r_data[4531] <= r_data[4530];
                
                r_data[4532] <= r_data[4531];
                
                r_data[4533] <= r_data[4532];
                
                r_data[4534] <= r_data[4533];
                
                r_data[4535] <= r_data[4534];
                
                r_data[4536] <= r_data[4535];
                
                r_data[4537] <= r_data[4536];
                
                r_data[4538] <= r_data[4537];
                
                r_data[4539] <= r_data[4538];
                
                r_data[4540] <= r_data[4539];
                
                r_data[4541] <= r_data[4540];
                
                r_data[4542] <= r_data[4541];
                
                r_data[4543] <= r_data[4542];
                
                r_data[4544] <= r_data[4543];
                
                r_data[4545] <= r_data[4544];
                
                r_data[4546] <= r_data[4545];
                
                r_data[4547] <= r_data[4546];
                
                r_data[4548] <= r_data[4547];
                
                r_data[4549] <= r_data[4548];
                
                r_data[4550] <= r_data[4549];
                
                r_data[4551] <= r_data[4550];
                
                r_data[4552] <= r_data[4551];
                
                r_data[4553] <= r_data[4552];
                
                r_data[4554] <= r_data[4553];
                
                r_data[4555] <= r_data[4554];
                
                r_data[4556] <= r_data[4555];
                
                r_data[4557] <= r_data[4556];
                
                r_data[4558] <= r_data[4557];
                
                r_data[4559] <= r_data[4558];
                
                r_data[4560] <= r_data[4559];
                
                r_data[4561] <= r_data[4560];
                
                r_data[4562] <= r_data[4561];
                
                r_data[4563] <= r_data[4562];
                
                r_data[4564] <= r_data[4563];
                
                r_data[4565] <= r_data[4564];
                
                r_data[4566] <= r_data[4565];
                
                r_data[4567] <= r_data[4566];
                
                r_data[4568] <= r_data[4567];
                
                r_data[4569] <= r_data[4568];
                
                r_data[4570] <= r_data[4569];
                
                r_data[4571] <= r_data[4570];
                
                r_data[4572] <= r_data[4571];
                
                r_data[4573] <= r_data[4572];
                
                r_data[4574] <= r_data[4573];
                
                r_data[4575] <= r_data[4574];
                
                r_data[4576] <= r_data[4575];
                
                r_data[4577] <= r_data[4576];
                
                r_data[4578] <= r_data[4577];
                
                r_data[4579] <= r_data[4578];
                
                r_data[4580] <= r_data[4579];
                
                r_data[4581] <= r_data[4580];
                
                r_data[4582] <= r_data[4581];
                
                r_data[4583] <= r_data[4582];
                
                r_data[4584] <= r_data[4583];
                
                r_data[4585] <= r_data[4584];
                
                r_data[4586] <= r_data[4585];
                
                r_data[4587] <= r_data[4586];
                
                r_data[4588] <= r_data[4587];
                
                r_data[4589] <= r_data[4588];
                
                r_data[4590] <= r_data[4589];
                
                r_data[4591] <= r_data[4590];
                
                r_data[4592] <= r_data[4591];
                
                r_data[4593] <= r_data[4592];
                
                r_data[4594] <= r_data[4593];
                
                r_data[4595] <= r_data[4594];
                
                r_data[4596] <= r_data[4595];
                
                r_data[4597] <= r_data[4596];
                
                r_data[4598] <= r_data[4597];
                
                r_data[4599] <= r_data[4598];
                
                r_data[4600] <= r_data[4599];
                
                r_data[4601] <= r_data[4600];
                
                r_data[4602] <= r_data[4601];
                
                r_data[4603] <= r_data[4602];
                
                r_data[4604] <= r_data[4603];
                
                r_data[4605] <= r_data[4604];
                
                r_data[4606] <= r_data[4605];
                
                r_data[4607] <= r_data[4606];
                
                r_data[4608] <= r_data[4607];
                
                r_data[4609] <= r_data[4608];
                
                r_data[4610] <= r_data[4609];
                
                r_data[4611] <= r_data[4610];
                
                r_data[4612] <= r_data[4611];
                
                r_data[4613] <= r_data[4612];
                
                r_data[4614] <= r_data[4613];
                
                r_data[4615] <= r_data[4614];
                
                r_data[4616] <= r_data[4615];
                
                r_data[4617] <= r_data[4616];
                
                r_data[4618] <= r_data[4617];
                
                r_data[4619] <= r_data[4618];
                
                r_data[4620] <= r_data[4619];
                
                r_data[4621] <= r_data[4620];
                
                r_data[4622] <= r_data[4621];
                
                r_data[4623] <= r_data[4622];
                
                r_data[4624] <= r_data[4623];
                
                r_data[4625] <= r_data[4624];
                
                r_data[4626] <= r_data[4625];
                
                r_data[4627] <= r_data[4626];
                
                r_data[4628] <= r_data[4627];
                
                r_data[4629] <= r_data[4628];
                
                r_data[4630] <= r_data[4629];
                
                r_data[4631] <= r_data[4630];
                
                r_data[4632] <= r_data[4631];
                
                r_data[4633] <= r_data[4632];
                
                r_data[4634] <= r_data[4633];
                
                r_data[4635] <= r_data[4634];
                
                r_data[4636] <= r_data[4635];
                
                r_data[4637] <= r_data[4636];
                
                r_data[4638] <= r_data[4637];
                
                r_data[4639] <= r_data[4638];
                
                r_data[4640] <= r_data[4639];
                
                r_data[4641] <= r_data[4640];
                
                r_data[4642] <= r_data[4641];
                
                r_data[4643] <= r_data[4642];
                
                r_data[4644] <= r_data[4643];
                
                r_data[4645] <= r_data[4644];
                
                r_data[4646] <= r_data[4645];
                
                r_data[4647] <= r_data[4646];
                
                r_data[4648] <= r_data[4647];
                
                r_data[4649] <= r_data[4648];
                
                r_data[4650] <= r_data[4649];
                
                r_data[4651] <= r_data[4650];
                
                r_data[4652] <= r_data[4651];
                
                r_data[4653] <= r_data[4652];
                
                r_data[4654] <= r_data[4653];
                
                r_data[4655] <= r_data[4654];
                
                r_data[4656] <= r_data[4655];
                
                r_data[4657] <= r_data[4656];
                
                r_data[4658] <= r_data[4657];
                
                r_data[4659] <= r_data[4658];
                
                r_data[4660] <= r_data[4659];
                
                r_data[4661] <= r_data[4660];
                
                r_data[4662] <= r_data[4661];
                
                r_data[4663] <= r_data[4662];
                
                r_data[4664] <= r_data[4663];
                
                r_data[4665] <= r_data[4664];
                
                r_data[4666] <= r_data[4665];
                
                r_data[4667] <= r_data[4666];
                
                r_data[4668] <= r_data[4667];
                
                r_data[4669] <= r_data[4668];
                
                r_data[4670] <= r_data[4669];
                
                r_data[4671] <= r_data[4670];
                
                r_data[4672] <= r_data[4671];
                
                r_data[4673] <= r_data[4672];
                
                r_data[4674] <= r_data[4673];
                
                r_data[4675] <= r_data[4674];
                
                r_data[4676] <= r_data[4675];
                
                r_data[4677] <= r_data[4676];
                
                r_data[4678] <= r_data[4677];
                
                r_data[4679] <= r_data[4678];
                
                r_data[4680] <= r_data[4679];
                
                r_data[4681] <= r_data[4680];
                
                r_data[4682] <= r_data[4681];
                
                r_data[4683] <= r_data[4682];
                
                r_data[4684] <= r_data[4683];
                
                r_data[4685] <= r_data[4684];
                
                r_data[4686] <= r_data[4685];
                
                r_data[4687] <= r_data[4686];
                
                r_data[4688] <= r_data[4687];
                
                r_data[4689] <= r_data[4688];
                
                r_data[4690] <= r_data[4689];
                
                r_data[4691] <= r_data[4690];
                
                r_data[4692] <= r_data[4691];
                
                r_data[4693] <= r_data[4692];
                
                r_data[4694] <= r_data[4693];
                
                r_data[4695] <= r_data[4694];
                
                r_data[4696] <= r_data[4695];
                
                r_data[4697] <= r_data[4696];
                
                r_data[4698] <= r_data[4697];
                
                r_data[4699] <= r_data[4698];
                
                r_data[4700] <= r_data[4699];
                
                r_data[4701] <= r_data[4700];
                
                r_data[4702] <= r_data[4701];
                
                r_data[4703] <= r_data[4702];
                
                r_data[4704] <= r_data[4703];
                
                r_data[4705] <= r_data[4704];
                
                r_data[4706] <= r_data[4705];
                
                r_data[4707] <= r_data[4706];
                
                r_data[4708] <= r_data[4707];
                
                r_data[4709] <= r_data[4708];
                
                r_data[4710] <= r_data[4709];
                
                r_data[4711] <= r_data[4710];
                
                r_data[4712] <= r_data[4711];
                
                r_data[4713] <= r_data[4712];
                
                r_data[4714] <= r_data[4713];
                
                r_data[4715] <= r_data[4714];
                
                r_data[4716] <= r_data[4715];
                
                r_data[4717] <= r_data[4716];
                
                r_data[4718] <= r_data[4717];
                
                r_data[4719] <= r_data[4718];
                
                r_data[4720] <= r_data[4719];
                
                r_data[4721] <= r_data[4720];
                
                r_data[4722] <= r_data[4721];
                
                r_data[4723] <= r_data[4722];
                
                r_data[4724] <= r_data[4723];
                
                r_data[4725] <= r_data[4724];
                
                r_data[4726] <= r_data[4725];
                
                r_data[4727] <= r_data[4726];
                
                r_data[4728] <= r_data[4727];
                
                r_data[4729] <= r_data[4728];
                
                r_data[4730] <= r_data[4729];
                
                r_data[4731] <= r_data[4730];
                
                r_data[4732] <= r_data[4731];
                
                r_data[4733] <= r_data[4732];
                
                r_data[4734] <= r_data[4733];
                
                r_data[4735] <= r_data[4734];
                
                r_data[4736] <= r_data[4735];
                
                r_data[4737] <= r_data[4736];
                
                r_data[4738] <= r_data[4737];
                
                r_data[4739] <= r_data[4738];
                
                r_data[4740] <= r_data[4739];
                
                r_data[4741] <= r_data[4740];
                
                r_data[4742] <= r_data[4741];
                
                r_data[4743] <= r_data[4742];
                
                r_data[4744] <= r_data[4743];
                
                r_data[4745] <= r_data[4744];
                
                r_data[4746] <= r_data[4745];
                
                r_data[4747] <= r_data[4746];
                
                r_data[4748] <= r_data[4747];
                
                r_data[4749] <= r_data[4748];
                
                r_data[4750] <= r_data[4749];
                
                r_data[4751] <= r_data[4750];
                
                r_data[4752] <= r_data[4751];
                
                r_data[4753] <= r_data[4752];
                
                r_data[4754] <= r_data[4753];
                
                r_data[4755] <= r_data[4754];
                
                r_data[4756] <= r_data[4755];
                
                r_data[4757] <= r_data[4756];
                
                r_data[4758] <= r_data[4757];
                
                r_data[4759] <= r_data[4758];
                
                r_data[4760] <= r_data[4759];
                
                r_data[4761] <= r_data[4760];
                
                r_data[4762] <= r_data[4761];
                
                r_data[4763] <= r_data[4762];
                
                r_data[4764] <= r_data[4763];
                
                r_data[4765] <= r_data[4764];
                
                r_data[4766] <= r_data[4765];
                
                r_data[4767] <= r_data[4766];
                
                r_data[4768] <= r_data[4767];
                
                r_data[4769] <= r_data[4768];
                
                r_data[4770] <= r_data[4769];
                
                r_data[4771] <= r_data[4770];
                
                r_data[4772] <= r_data[4771];
                
                r_data[4773] <= r_data[4772];
                
                r_data[4774] <= r_data[4773];
                
                r_data[4775] <= r_data[4774];
                
                r_data[4776] <= r_data[4775];
                
                r_data[4777] <= r_data[4776];
                
                r_data[4778] <= r_data[4777];
                
                r_data[4779] <= r_data[4778];
                
                r_data[4780] <= r_data[4779];
                
                r_data[4781] <= r_data[4780];
                
                r_data[4782] <= r_data[4781];
                
                r_data[4783] <= r_data[4782];
                
                r_data[4784] <= r_data[4783];
                
                r_data[4785] <= r_data[4784];
                
                r_data[4786] <= r_data[4785];
                
                r_data[4787] <= r_data[4786];
                
                r_data[4788] <= r_data[4787];
                
                r_data[4789] <= r_data[4788];
                
                r_data[4790] <= r_data[4789];
                
                r_data[4791] <= r_data[4790];
                
                r_data[4792] <= r_data[4791];
                
                r_data[4793] <= r_data[4792];
                
                r_data[4794] <= r_data[4793];
                
                r_data[4795] <= r_data[4794];
                
                r_data[4796] <= r_data[4795];
                
                r_data[4797] <= r_data[4796];
                
                r_data[4798] <= r_data[4797];
                
                r_data[4799] <= r_data[4798];
                
                r_data[4800] <= r_data[4799];
                
                r_data[4801] <= r_data[4800];
                
                r_data[4802] <= r_data[4801];
                
                r_data[4803] <= r_data[4802];
                
                r_data[4804] <= r_data[4803];
                
                r_data[4805] <= r_data[4804];
                
                r_data[4806] <= r_data[4805];
                
                r_data[4807] <= r_data[4806];
                
                r_data[4808] <= r_data[4807];
                
                r_data[4809] <= r_data[4808];
                
                r_data[4810] <= r_data[4809];
                
                r_data[4811] <= r_data[4810];
                
                r_data[4812] <= r_data[4811];
                
                r_data[4813] <= r_data[4812];
                
                r_data[4814] <= r_data[4813];
                
                r_data[4815] <= r_data[4814];
                
                r_data[4816] <= r_data[4815];
                
                r_data[4817] <= r_data[4816];
                
                r_data[4818] <= r_data[4817];
                
                r_data[4819] <= r_data[4818];
                
                r_data[4820] <= r_data[4819];
                
                r_data[4821] <= r_data[4820];
                
                r_data[4822] <= r_data[4821];
                
                r_data[4823] <= r_data[4822];
                
                r_data[4824] <= r_data[4823];
                
                r_data[4825] <= r_data[4824];
                
                r_data[4826] <= r_data[4825];
                
                r_data[4827] <= r_data[4826];
                
                r_data[4828] <= r_data[4827];
                
                r_data[4829] <= r_data[4828];
                
                r_data[4830] <= r_data[4829];
                
                r_data[4831] <= r_data[4830];
                
                r_data[4832] <= r_data[4831];
                
                r_data[4833] <= r_data[4832];
                
                r_data[4834] <= r_data[4833];
                
                r_data[4835] <= r_data[4834];
                
                r_data[4836] <= r_data[4835];
                
                r_data[4837] <= r_data[4836];
                
                r_data[4838] <= r_data[4837];
                
                r_data[4839] <= r_data[4838];
                
                r_data[4840] <= r_data[4839];
                
                r_data[4841] <= r_data[4840];
                
                r_data[4842] <= r_data[4841];
                
                r_data[4843] <= r_data[4842];
                
                r_data[4844] <= r_data[4843];
                
                r_data[4845] <= r_data[4844];
                
                r_data[4846] <= r_data[4845];
                
                r_data[4847] <= r_data[4846];
                
                r_data[4848] <= r_data[4847];
                
                r_data[4849] <= r_data[4848];
                
                r_data[4850] <= r_data[4849];
                
                r_data[4851] <= r_data[4850];
                
                r_data[4852] <= r_data[4851];
                
                r_data[4853] <= r_data[4852];
                
                r_data[4854] <= r_data[4853];
                
                r_data[4855] <= r_data[4854];
                
                r_data[4856] <= r_data[4855];
                
                r_data[4857] <= r_data[4856];
                
                r_data[4858] <= r_data[4857];
                
                r_data[4859] <= r_data[4858];
                
                r_data[4860] <= r_data[4859];
                
                r_data[4861] <= r_data[4860];
                
                r_data[4862] <= r_data[4861];
                
                r_data[4863] <= r_data[4862];
                
                r_data[4864] <= r_data[4863];
                
                r_data[4865] <= r_data[4864];
                
                r_data[4866] <= r_data[4865];
                
                r_data[4867] <= r_data[4866];
                
                r_data[4868] <= r_data[4867];
                
                r_data[4869] <= r_data[4868];
                
                r_data[4870] <= r_data[4869];
                
                r_data[4871] <= r_data[4870];
                
                r_data[4872] <= r_data[4871];
                
                r_data[4873] <= r_data[4872];
                
                r_data[4874] <= r_data[4873];
                
                r_data[4875] <= r_data[4874];
                
                r_data[4876] <= r_data[4875];
                
                r_data[4877] <= r_data[4876];
                
                r_data[4878] <= r_data[4877];
                
                r_data[4879] <= r_data[4878];
                
                r_data[4880] <= r_data[4879];
                
                r_data[4881] <= r_data[4880];
                
                r_data[4882] <= r_data[4881];
                
                r_data[4883] <= r_data[4882];
                
                r_data[4884] <= r_data[4883];
                
                r_data[4885] <= r_data[4884];
                
                r_data[4886] <= r_data[4885];
                
                r_data[4887] <= r_data[4886];
                
                r_data[4888] <= r_data[4887];
                
                r_data[4889] <= r_data[4888];
                
                r_data[4890] <= r_data[4889];
                
                r_data[4891] <= r_data[4890];
                
                r_data[4892] <= r_data[4891];
                
                r_data[4893] <= r_data[4892];
                
                r_data[4894] <= r_data[4893];
                
                r_data[4895] <= r_data[4894];
                
                r_data[4896] <= r_data[4895];
                
                r_data[4897] <= r_data[4896];
                
                r_data[4898] <= r_data[4897];
                
                r_data[4899] <= r_data[4898];
                
                r_data[4900] <= r_data[4899];
                
                r_data[4901] <= r_data[4900];
                
                r_data[4902] <= r_data[4901];
                
                r_data[4903] <= r_data[4902];
                
                r_data[4904] <= r_data[4903];
                
                r_data[4905] <= r_data[4904];
                
                r_data[4906] <= r_data[4905];
                
                r_data[4907] <= r_data[4906];
                
                r_data[4908] <= r_data[4907];
                
                r_data[4909] <= r_data[4908];
                
                r_data[4910] <= r_data[4909];
                
                r_data[4911] <= r_data[4910];
                
                r_data[4912] <= r_data[4911];
                
                r_data[4913] <= r_data[4912];
                
                r_data[4914] <= r_data[4913];
                
                r_data[4915] <= r_data[4914];
                
                r_data[4916] <= r_data[4915];
                
                r_data[4917] <= r_data[4916];
                
                r_data[4918] <= r_data[4917];
                
                r_data[4919] <= r_data[4918];
                
                r_data[4920] <= r_data[4919];
                
                r_data[4921] <= r_data[4920];
                
                r_data[4922] <= r_data[4921];
                
                r_data[4923] <= r_data[4922];
                
                r_data[4924] <= r_data[4923];
                
                r_data[4925] <= r_data[4924];
                
                r_data[4926] <= r_data[4925];
                
                r_data[4927] <= r_data[4926];
                
                r_data[4928] <= r_data[4927];
                
                r_data[4929] <= r_data[4928];
                
                r_data[4930] <= r_data[4929];
                
                r_data[4931] <= r_data[4930];
                
                r_data[4932] <= r_data[4931];
                
                r_data[4933] <= r_data[4932];
                
                r_data[4934] <= r_data[4933];
                
                r_data[4935] <= r_data[4934];
                
                r_data[4936] <= r_data[4935];
                
                r_data[4937] <= r_data[4936];
                
                r_data[4938] <= r_data[4937];
                
                r_data[4939] <= r_data[4938];
                
                r_data[4940] <= r_data[4939];
                
                r_data[4941] <= r_data[4940];
                
                r_data[4942] <= r_data[4941];
                
                r_data[4943] <= r_data[4942];
                
                r_data[4944] <= r_data[4943];
                
                r_data[4945] <= r_data[4944];
                
                r_data[4946] <= r_data[4945];
                
                r_data[4947] <= r_data[4946];
                
                r_data[4948] <= r_data[4947];
                
                r_data[4949] <= r_data[4948];
                
                r_data[4950] <= r_data[4949];
                
                r_data[4951] <= r_data[4950];
                
                r_data[4952] <= r_data[4951];
                
                r_data[4953] <= r_data[4952];
                
                r_data[4954] <= r_data[4953];
                
                r_data[4955] <= r_data[4954];
                
                r_data[4956] <= r_data[4955];
                
                r_data[4957] <= r_data[4956];
                
                r_data[4958] <= r_data[4957];
                
                r_data[4959] <= r_data[4958];
                
                r_data[4960] <= r_data[4959];
                
                r_data[4961] <= r_data[4960];
                
                r_data[4962] <= r_data[4961];
                
                r_data[4963] <= r_data[4962];
                
                r_data[4964] <= r_data[4963];
                
                r_data[4965] <= r_data[4964];
                
                r_data[4966] <= r_data[4965];
                
                r_data[4967] <= r_data[4966];
                
                r_data[4968] <= r_data[4967];
                
                r_data[4969] <= r_data[4968];
                
                r_data[4970] <= r_data[4969];
                
                r_data[4971] <= r_data[4970];
                
                r_data[4972] <= r_data[4971];
                
                r_data[4973] <= r_data[4972];
                
                r_data[4974] <= r_data[4973];
                
                r_data[4975] <= r_data[4974];
                
                r_data[4976] <= r_data[4975];
                
                r_data[4977] <= r_data[4976];
                
                r_data[4978] <= r_data[4977];
                
                r_data[4979] <= r_data[4978];
                
                r_data[4980] <= r_data[4979];
                
                r_data[4981] <= r_data[4980];
                
                r_data[4982] <= r_data[4981];
                
                r_data[4983] <= r_data[4982];
                
                r_data[4984] <= r_data[4983];
                
                r_data[4985] <= r_data[4984];
                
                r_data[4986] <= r_data[4985];
                
                r_data[4987] <= r_data[4986];
                
                r_data[4988] <= r_data[4987];
                
                r_data[4989] <= r_data[4988];
                
                r_data[4990] <= r_data[4989];
                
                r_data[4991] <= r_data[4990];
                
                r_data[4992] <= r_data[4991];
                
                r_data[4993] <= r_data[4992];
                
                r_data[4994] <= r_data[4993];
                
                r_data[4995] <= r_data[4994];
                
                r_data[4996] <= r_data[4995];
                
                r_data[4997] <= r_data[4996];
                
                r_data[4998] <= r_data[4997];
                
                r_data[4999] <= r_data[4998];
                
                r_data[5000] <= r_data[4999];
                
                r_data[5001] <= r_data[5000];
                
                r_data[5002] <= r_data[5001];
                
                r_data[5003] <= r_data[5002];
                
                r_data[5004] <= r_data[5003];
                
                r_data[5005] <= r_data[5004];
                
                r_data[5006] <= r_data[5005];
                
                r_data[5007] <= r_data[5006];
                
                r_data[5008] <= r_data[5007];
                
                r_data[5009] <= r_data[5008];
                
                r_data[5010] <= r_data[5009];
                
                r_data[5011] <= r_data[5010];
                
                r_data[5012] <= r_data[5011];
                
                r_data[5013] <= r_data[5012];
                
                r_data[5014] <= r_data[5013];
                
                r_data[5015] <= r_data[5014];
                
                r_data[5016] <= r_data[5015];
                
                r_data[5017] <= r_data[5016];
                
                r_data[5018] <= r_data[5017];
                
                r_data[5019] <= r_data[5018];
                
                r_data[5020] <= r_data[5019];
                
                r_data[5021] <= r_data[5020];
                
                r_data[5022] <= r_data[5021];
                
                r_data[5023] <= r_data[5022];
                
                r_data[5024] <= r_data[5023];
                
                r_data[5025] <= r_data[5024];
                
                r_data[5026] <= r_data[5025];
                
                r_data[5027] <= r_data[5026];
                
                r_data[5028] <= r_data[5027];
                
                r_data[5029] <= r_data[5028];
                
                r_data[5030] <= r_data[5029];
                
                r_data[5031] <= r_data[5030];
                
                r_data[5032] <= r_data[5031];
                
                r_data[5033] <= r_data[5032];
                
                r_data[5034] <= r_data[5033];
                
                r_data[5035] <= r_data[5034];
                
                r_data[5036] <= r_data[5035];
                
                r_data[5037] <= r_data[5036];
                
                r_data[5038] <= r_data[5037];
                
                r_data[5039] <= r_data[5038];
                
                r_data[5040] <= r_data[5039];
                
                r_data[5041] <= r_data[5040];
                
                r_data[5042] <= r_data[5041];
                
                r_data[5043] <= r_data[5042];
                
                r_data[5044] <= r_data[5043];
                
                r_data[5045] <= r_data[5044];
                
                r_data[5046] <= r_data[5045];
                
                r_data[5047] <= r_data[5046];
                
                r_data[5048] <= r_data[5047];
                
                r_data[5049] <= r_data[5048];
                
                r_data[5050] <= r_data[5049];
                
                r_data[5051] <= r_data[5050];
                
                r_data[5052] <= r_data[5051];
                
                r_data[5053] <= r_data[5052];
                
                r_data[5054] <= r_data[5053];
                
                r_data[5055] <= r_data[5054];
                
                r_data[5056] <= r_data[5055];
                
                r_data[5057] <= r_data[5056];
                
                r_data[5058] <= r_data[5057];
                
                r_data[5059] <= r_data[5058];
                
                r_data[5060] <= r_data[5059];
                
                r_data[5061] <= r_data[5060];
                
                r_data[5062] <= r_data[5061];
                
                r_data[5063] <= r_data[5062];
                
                r_data[5064] <= r_data[5063];
                
                r_data[5065] <= r_data[5064];
                
                r_data[5066] <= r_data[5065];
                
                r_data[5067] <= r_data[5066];
                
                r_data[5068] <= r_data[5067];
                
                r_data[5069] <= r_data[5068];
                
                r_data[5070] <= r_data[5069];
                
                r_data[5071] <= r_data[5070];
                
                r_data[5072] <= r_data[5071];
                
                r_data[5073] <= r_data[5072];
                
                r_data[5074] <= r_data[5073];
                
                r_data[5075] <= r_data[5074];
                
                r_data[5076] <= r_data[5075];
                
                r_data[5077] <= r_data[5076];
                
                r_data[5078] <= r_data[5077];
                
                r_data[5079] <= r_data[5078];
                
                r_data[5080] <= r_data[5079];
                
                r_data[5081] <= r_data[5080];
                
                r_data[5082] <= r_data[5081];
                
                r_data[5083] <= r_data[5082];
                
                r_data[5084] <= r_data[5083];
                
                r_data[5085] <= r_data[5084];
                
                r_data[5086] <= r_data[5085];
                
                r_data[5087] <= r_data[5086];
                
                r_data[5088] <= r_data[5087];
                
                r_data[5089] <= r_data[5088];
                
                r_data[5090] <= r_data[5089];
                
                r_data[5091] <= r_data[5090];
                
                r_data[5092] <= r_data[5091];
                
                r_data[5093] <= r_data[5092];
                
                r_data[5094] <= r_data[5093];
                
                r_data[5095] <= r_data[5094];
                
                r_data[5096] <= r_data[5095];
                
                r_data[5097] <= r_data[5096];
                
                r_data[5098] <= r_data[5097];
                
                r_data[5099] <= r_data[5098];
                
                r_data[5100] <= r_data[5099];
                
                r_data[5101] <= r_data[5100];
                
                r_data[5102] <= r_data[5101];
                
                r_data[5103] <= r_data[5102];
                
                r_data[5104] <= r_data[5103];
                
                r_data[5105] <= r_data[5104];
                
                r_data[5106] <= r_data[5105];
                
                r_data[5107] <= r_data[5106];
                
                r_data[5108] <= r_data[5107];
                
                r_data[5109] <= r_data[5108];
                
                r_data[5110] <= r_data[5109];
                
                r_data[5111] <= r_data[5110];
                
                r_data[5112] <= r_data[5111];
                
                r_data[5113] <= r_data[5112];
                
                r_data[5114] <= r_data[5113];
                
                r_data[5115] <= r_data[5114];
                
                r_data[5116] <= r_data[5115];
                
                r_data[5117] <= r_data[5116];
                
                r_data[5118] <= r_data[5117];
                
                r_data[5119] <= r_data[5118];
                
                r_data[5120] <= r_data[5119];
                
                r_data[5121] <= r_data[5120];
                
                r_data[5122] <= r_data[5121];
                
                r_data[5123] <= r_data[5122];
                
                r_data[5124] <= r_data[5123];
                
                r_data[5125] <= r_data[5124];
                
                r_data[5126] <= r_data[5125];
                
                r_data[5127] <= r_data[5126];
                
                r_data[5128] <= r_data[5127];
                
                r_data[5129] <= r_data[5128];
                
                r_data[5130] <= r_data[5129];
                
                r_data[5131] <= r_data[5130];
                
                r_data[5132] <= r_data[5131];
                
                r_data[5133] <= r_data[5132];
                
                r_data[5134] <= r_data[5133];
                
                r_data[5135] <= r_data[5134];
                
                r_data[5136] <= r_data[5135];
                
                r_data[5137] <= r_data[5136];
                
                r_data[5138] <= r_data[5137];
                
                r_data[5139] <= r_data[5138];
                
                r_data[5140] <= r_data[5139];
                
                r_data[5141] <= r_data[5140];
                
                r_data[5142] <= r_data[5141];
                
                r_data[5143] <= r_data[5142];
                
                r_data[5144] <= r_data[5143];
                
                r_data[5145] <= r_data[5144];
                
                r_data[5146] <= r_data[5145];
                
                r_data[5147] <= r_data[5146];
                
                r_data[5148] <= r_data[5147];
                
                r_data[5149] <= r_data[5148];
                
                r_data[5150] <= r_data[5149];
                
                r_data[5151] <= r_data[5150];
                
                r_data[5152] <= r_data[5151];
                
                r_data[5153] <= r_data[5152];
                
                r_data[5154] <= r_data[5153];
                
                r_data[5155] <= r_data[5154];
                
                r_data[5156] <= r_data[5155];
                
                r_data[5157] <= r_data[5156];
                
                r_data[5158] <= r_data[5157];
                
                r_data[5159] <= r_data[5158];
                
                r_data[5160] <= r_data[5159];
                
                r_data[5161] <= r_data[5160];
                
                r_data[5162] <= r_data[5161];
                
                r_data[5163] <= r_data[5162];
                
                r_data[5164] <= r_data[5163];
                
                r_data[5165] <= r_data[5164];
                
                r_data[5166] <= r_data[5165];
                
                r_data[5167] <= r_data[5166];
                
                r_data[5168] <= r_data[5167];
                
                r_data[5169] <= r_data[5168];
                
                r_data[5170] <= r_data[5169];
                
                r_data[5171] <= r_data[5170];
                
                r_data[5172] <= r_data[5171];
                
                r_data[5173] <= r_data[5172];
                
                r_data[5174] <= r_data[5173];
                
                r_data[5175] <= r_data[5174];
                
                r_data[5176] <= r_data[5175];
                
                r_data[5177] <= r_data[5176];
                
                r_data[5178] <= r_data[5177];
                
                r_data[5179] <= r_data[5178];
                
                r_data[5180] <= r_data[5179];
                
                r_data[5181] <= r_data[5180];
                
                r_data[5182] <= r_data[5181];
                
                r_data[5183] <= r_data[5182];
                
                r_data[5184] <= r_data[5183];
                
                r_data[5185] <= r_data[5184];
                
                r_data[5186] <= r_data[5185];
                
                r_data[5187] <= r_data[5186];
                
                r_data[5188] <= r_data[5187];
                
                r_data[5189] <= r_data[5188];
                
                r_data[5190] <= r_data[5189];
                
                r_data[5191] <= r_data[5190];
                
                r_data[5192] <= r_data[5191];
                
                r_data[5193] <= r_data[5192];
                
                r_data[5194] <= r_data[5193];
                
                r_data[5195] <= r_data[5194];
                
                r_data[5196] <= r_data[5195];
                
                r_data[5197] <= r_data[5196];
                
                r_data[5198] <= r_data[5197];
                
                r_data[5199] <= r_data[5198];
                
                r_data[5200] <= r_data[5199];
                
                r_data[5201] <= r_data[5200];
                
                r_data[5202] <= r_data[5201];
                
                r_data[5203] <= r_data[5202];
                
                r_data[5204] <= r_data[5203];
                
                r_data[5205] <= r_data[5204];
                
                r_data[5206] <= r_data[5205];
                
                r_data[5207] <= r_data[5206];
                
                r_data[5208] <= r_data[5207];
                
                r_data[5209] <= r_data[5208];
                
                r_data[5210] <= r_data[5209];
                
                r_data[5211] <= r_data[5210];
                
                r_data[5212] <= r_data[5211];
                
                r_data[5213] <= r_data[5212];
                
                r_data[5214] <= r_data[5213];
                
                r_data[5215] <= r_data[5214];
                
                r_data[5216] <= r_data[5215];
                
                r_data[5217] <= r_data[5216];
                
                r_data[5218] <= r_data[5217];
                
                r_data[5219] <= r_data[5218];
                
                r_data[5220] <= r_data[5219];
                
                r_data[5221] <= r_data[5220];
                
                r_data[5222] <= r_data[5221];
                
                r_data[5223] <= r_data[5222];
                
                r_data[5224] <= r_data[5223];
                
                r_data[5225] <= r_data[5224];
                
                r_data[5226] <= r_data[5225];
                
                r_data[5227] <= r_data[5226];
                
                r_data[5228] <= r_data[5227];
                
                r_data[5229] <= r_data[5228];
                
                r_data[5230] <= r_data[5229];
                
                r_data[5231] <= r_data[5230];
                
                r_data[5232] <= r_data[5231];
                
                r_data[5233] <= r_data[5232];
                
                r_data[5234] <= r_data[5233];
                
                r_data[5235] <= r_data[5234];
                
                r_data[5236] <= r_data[5235];
                
                r_data[5237] <= r_data[5236];
                
                r_data[5238] <= r_data[5237];
                
                r_data[5239] <= r_data[5238];
                
                r_data[5240] <= r_data[5239];
                
                r_data[5241] <= r_data[5240];
                
                r_data[5242] <= r_data[5241];
                
                r_data[5243] <= r_data[5242];
                
                r_data[5244] <= r_data[5243];
                
                r_data[5245] <= r_data[5244];
                
                r_data[5246] <= r_data[5245];
                
                r_data[5247] <= r_data[5246];
                
                r_data[5248] <= r_data[5247];
                
                r_data[5249] <= r_data[5248];
                
                r_data[5250] <= r_data[5249];
                
                r_data[5251] <= r_data[5250];
                
                r_data[5252] <= r_data[5251];
                
                r_data[5253] <= r_data[5252];
                
                r_data[5254] <= r_data[5253];
                
                r_data[5255] <= r_data[5254];
                
                r_data[5256] <= r_data[5255];
                
                r_data[5257] <= r_data[5256];
                
                r_data[5258] <= r_data[5257];
                
                r_data[5259] <= r_data[5258];
                
                r_data[5260] <= r_data[5259];
                
                r_data[5261] <= r_data[5260];
                
                r_data[5262] <= r_data[5261];
                
                r_data[5263] <= r_data[5262];
                
                r_data[5264] <= r_data[5263];
                
                r_data[5265] <= r_data[5264];
                
                r_data[5266] <= r_data[5265];
                
                r_data[5267] <= r_data[5266];
                
                r_data[5268] <= r_data[5267];
                
                r_data[5269] <= r_data[5268];
                
                r_data[5270] <= r_data[5269];
                
                r_data[5271] <= r_data[5270];
                
                r_data[5272] <= r_data[5271];
                
                r_data[5273] <= r_data[5272];
                
                r_data[5274] <= r_data[5273];
                
                r_data[5275] <= r_data[5274];
                
                r_data[5276] <= r_data[5275];
                
                r_data[5277] <= r_data[5276];
                
                r_data[5278] <= r_data[5277];
                
                r_data[5279] <= r_data[5278];
                
                r_data[5280] <= r_data[5279];
                
                r_data[5281] <= r_data[5280];
                
                r_data[5282] <= r_data[5281];
                
                r_data[5283] <= r_data[5282];
                
                r_data[5284] <= r_data[5283];
                
                r_data[5285] <= r_data[5284];
                
                r_data[5286] <= r_data[5285];
                
                r_data[5287] <= r_data[5286];
                
                r_data[5288] <= r_data[5287];
                
                r_data[5289] <= r_data[5288];
                
                r_data[5290] <= r_data[5289];
                
                r_data[5291] <= r_data[5290];
                
                r_data[5292] <= r_data[5291];
                
                r_data[5293] <= r_data[5292];
                
                r_data[5294] <= r_data[5293];
                
                r_data[5295] <= r_data[5294];
                
                r_data[5296] <= r_data[5295];
                
                r_data[5297] <= r_data[5296];
                
                r_data[5298] <= r_data[5297];
                
                r_data[5299] <= r_data[5298];
                
                r_data[5300] <= r_data[5299];
                
                r_data[5301] <= r_data[5300];
                
                r_data[5302] <= r_data[5301];
                
                r_data[5303] <= r_data[5302];
                
                r_data[5304] <= r_data[5303];
                
                r_data[5305] <= r_data[5304];
                
                r_data[5306] <= r_data[5305];
                
                r_data[5307] <= r_data[5306];
                
                r_data[5308] <= r_data[5307];
                
                r_data[5309] <= r_data[5308];
                
                r_data[5310] <= r_data[5309];
                
                r_data[5311] <= r_data[5310];
                
                r_data[5312] <= r_data[5311];
                
                r_data[5313] <= r_data[5312];
                
                r_data[5314] <= r_data[5313];
                
                r_data[5315] <= r_data[5314];
                
                r_data[5316] <= r_data[5315];
                
                r_data[5317] <= r_data[5316];
                
                r_data[5318] <= r_data[5317];
                
                r_data[5319] <= r_data[5318];
                
                r_data[5320] <= r_data[5319];
                
                r_data[5321] <= r_data[5320];
                
                r_data[5322] <= r_data[5321];
                
                r_data[5323] <= r_data[5322];
                
                r_data[5324] <= r_data[5323];
                
                r_data[5325] <= r_data[5324];
                
                r_data[5326] <= r_data[5325];
                
                r_data[5327] <= r_data[5326];
                
                r_data[5328] <= r_data[5327];
                
                r_data[5329] <= r_data[5328];
                
                r_data[5330] <= r_data[5329];
                
                r_data[5331] <= r_data[5330];
                
                r_data[5332] <= r_data[5331];
                
                r_data[5333] <= r_data[5332];
                
                r_data[5334] <= r_data[5333];
                
                r_data[5335] <= r_data[5334];
                
                r_data[5336] <= r_data[5335];
                
                r_data[5337] <= r_data[5336];
                
                r_data[5338] <= r_data[5337];
                
                r_data[5339] <= r_data[5338];
                
                r_data[5340] <= r_data[5339];
                
                r_data[5341] <= r_data[5340];
                
                r_data[5342] <= r_data[5341];
                
                r_data[5343] <= r_data[5342];
                
                r_data[5344] <= r_data[5343];
                
                r_data[5345] <= r_data[5344];
                
                r_data[5346] <= r_data[5345];
                
                r_data[5347] <= r_data[5346];
                
                r_data[5348] <= r_data[5347];
                
                r_data[5349] <= r_data[5348];
                
                r_data[5350] <= r_data[5349];
                
                r_data[5351] <= r_data[5350];
                
                r_data[5352] <= r_data[5351];
                
                r_data[5353] <= r_data[5352];
                
                r_data[5354] <= r_data[5353];
                
                r_data[5355] <= r_data[5354];
                
                r_data[5356] <= r_data[5355];
                
                r_data[5357] <= r_data[5356];
                
                r_data[5358] <= r_data[5357];
                
                r_data[5359] <= r_data[5358];
                
                r_data[5360] <= r_data[5359];
                
                r_data[5361] <= r_data[5360];
                
                r_data[5362] <= r_data[5361];
                
                r_data[5363] <= r_data[5362];
                
                r_data[5364] <= r_data[5363];
                
                r_data[5365] <= r_data[5364];
                
                r_data[5366] <= r_data[5365];
                
                r_data[5367] <= r_data[5366];
                
                r_data[5368] <= r_data[5367];
                
                r_data[5369] <= r_data[5368];
                
                r_data[5370] <= r_data[5369];
                
                r_data[5371] <= r_data[5370];
                
                r_data[5372] <= r_data[5371];
                
                r_data[5373] <= r_data[5372];
                
                r_data[5374] <= r_data[5373];
                
                r_data[5375] <= r_data[5374];
                
                r_data[5376] <= r_data[5375];
                
                r_data[5377] <= r_data[5376];
                
                r_data[5378] <= r_data[5377];
                
                r_data[5379] <= r_data[5378];
                
                r_data[5380] <= r_data[5379];
                
                r_data[5381] <= r_data[5380];
                
                r_data[5382] <= r_data[5381];
                
                r_data[5383] <= r_data[5382];
                
                r_data[5384] <= r_data[5383];
                
                r_data[5385] <= r_data[5384];
                
                r_data[5386] <= r_data[5385];
                
                r_data[5387] <= r_data[5386];
                
                r_data[5388] <= r_data[5387];
                
                r_data[5389] <= r_data[5388];
                
                r_data[5390] <= r_data[5389];
                
                r_data[5391] <= r_data[5390];
                
                r_data[5392] <= r_data[5391];
                
                r_data[5393] <= r_data[5392];
                
                r_data[5394] <= r_data[5393];
                
                r_data[5395] <= r_data[5394];
                
                r_data[5396] <= r_data[5395];
                
                r_data[5397] <= r_data[5396];
                
                r_data[5398] <= r_data[5397];
                
                r_data[5399] <= r_data[5398];
                
                r_data[5400] <= r_data[5399];
                
                r_data[5401] <= r_data[5400];
                
                r_data[5402] <= r_data[5401];
                
                r_data[5403] <= r_data[5402];
                
                r_data[5404] <= r_data[5403];
                
                r_data[5405] <= r_data[5404];
                
                r_data[5406] <= r_data[5405];
                
                r_data[5407] <= r_data[5406];
                
                r_data[5408] <= r_data[5407];
                
                r_data[5409] <= r_data[5408];
                
                r_data[5410] <= r_data[5409];
                
                r_data[5411] <= r_data[5410];
                
                r_data[5412] <= r_data[5411];
                
                r_data[5413] <= r_data[5412];
                
                r_data[5414] <= r_data[5413];
                
                r_data[5415] <= r_data[5414];
                
                r_data[5416] <= r_data[5415];
                
                r_data[5417] <= r_data[5416];
                
                r_data[5418] <= r_data[5417];
                
                r_data[5419] <= r_data[5418];
                
                r_data[5420] <= r_data[5419];
                
                r_data[5421] <= r_data[5420];
                
                r_data[5422] <= r_data[5421];
                
                r_data[5423] <= r_data[5422];
                
                r_data[5424] <= r_data[5423];
                
                r_data[5425] <= r_data[5424];
                
                r_data[5426] <= r_data[5425];
                
                r_data[5427] <= r_data[5426];
                
                r_data[5428] <= r_data[5427];
                
                r_data[5429] <= r_data[5428];
                
                r_data[5430] <= r_data[5429];
                
                r_data[5431] <= r_data[5430];
                
                r_data[5432] <= r_data[5431];
                
                r_data[5433] <= r_data[5432];
                
                r_data[5434] <= r_data[5433];
                
                r_data[5435] <= r_data[5434];
                
                r_data[5436] <= r_data[5435];
                
                r_data[5437] <= r_data[5436];
                
                r_data[5438] <= r_data[5437];
                
                r_data[5439] <= r_data[5438];
                
                r_data[5440] <= r_data[5439];
                
                r_data[5441] <= r_data[5440];
                
                r_data[5442] <= r_data[5441];
                
                r_data[5443] <= r_data[5442];
                
                r_data[5444] <= r_data[5443];
                
                r_data[5445] <= r_data[5444];
                
                r_data[5446] <= r_data[5445];
                
                r_data[5447] <= r_data[5446];
                
                r_data[5448] <= r_data[5447];
                
                r_data[5449] <= r_data[5448];
                
                r_data[5450] <= r_data[5449];
                
                r_data[5451] <= r_data[5450];
                
                r_data[5452] <= r_data[5451];
                
                r_data[5453] <= r_data[5452];
                
                r_data[5454] <= r_data[5453];
                
                r_data[5455] <= r_data[5454];
                
                r_data[5456] <= r_data[5455];
                
                r_data[5457] <= r_data[5456];
                
                r_data[5458] <= r_data[5457];
                
                r_data[5459] <= r_data[5458];
                
                r_data[5460] <= r_data[5459];
                
                r_data[5461] <= r_data[5460];
                
                r_data[5462] <= r_data[5461];
                
                r_data[5463] <= r_data[5462];
                
                r_data[5464] <= r_data[5463];
                
                r_data[5465] <= r_data[5464];
                
                r_data[5466] <= r_data[5465];
                
                r_data[5467] <= r_data[5466];
                
                r_data[5468] <= r_data[5467];
                
                r_data[5469] <= r_data[5468];
                
                r_data[5470] <= r_data[5469];
                
                r_data[5471] <= r_data[5470];
                
                r_data[5472] <= r_data[5471];
                
                r_data[5473] <= r_data[5472];
                
                r_data[5474] <= r_data[5473];
                
                r_data[5475] <= r_data[5474];
                
                r_data[5476] <= r_data[5475];
                
                r_data[5477] <= r_data[5476];
                
                r_data[5478] <= r_data[5477];
                
                r_data[5479] <= r_data[5478];
                
                r_data[5480] <= r_data[5479];
                
                r_data[5481] <= r_data[5480];
                
                r_data[5482] <= r_data[5481];
                
                r_data[5483] <= r_data[5482];
                
                r_data[5484] <= r_data[5483];
                
                r_data[5485] <= r_data[5484];
                
                r_data[5486] <= r_data[5485];
                
                r_data[5487] <= r_data[5486];
                
                r_data[5488] <= r_data[5487];
                
                r_data[5489] <= r_data[5488];
                
                r_data[5490] <= r_data[5489];
                
                r_data[5491] <= r_data[5490];
                
                r_data[5492] <= r_data[5491];
                
                r_data[5493] <= r_data[5492];
                
                r_data[5494] <= r_data[5493];
                
                r_data[5495] <= r_data[5494];
                
                r_data[5496] <= r_data[5495];
                
                r_data[5497] <= r_data[5496];
                
                r_data[5498] <= r_data[5497];
                
                r_data[5499] <= r_data[5498];
                
                r_data[5500] <= r_data[5499];
                
                r_data[5501] <= r_data[5500];
                
                r_data[5502] <= r_data[5501];
                
                r_data[5503] <= r_data[5502];
                
                r_data[5504] <= r_data[5503];
                
                r_data[5505] <= r_data[5504];
                
                r_data[5506] <= r_data[5505];
                
                r_data[5507] <= r_data[5506];
                
                r_data[5508] <= r_data[5507];
                
                r_data[5509] <= r_data[5508];
                
                r_data[5510] <= r_data[5509];
                
                r_data[5511] <= r_data[5510];
                
                r_data[5512] <= r_data[5511];
                
                r_data[5513] <= r_data[5512];
                
                r_data[5514] <= r_data[5513];
                
                r_data[5515] <= r_data[5514];
                
                r_data[5516] <= r_data[5515];
                
                r_data[5517] <= r_data[5516];
                
                r_data[5518] <= r_data[5517];
                
                r_data[5519] <= r_data[5518];
                
                r_data[5520] <= r_data[5519];
                
                r_data[5521] <= r_data[5520];
                
                r_data[5522] <= r_data[5521];
                
                r_data[5523] <= r_data[5522];
                
                r_data[5524] <= r_data[5523];
                
                r_data[5525] <= r_data[5524];
                
                r_data[5526] <= r_data[5525];
                
                r_data[5527] <= r_data[5526];
                
                r_data[5528] <= r_data[5527];
                
                r_data[5529] <= r_data[5528];
                
                r_data[5530] <= r_data[5529];
                
                r_data[5531] <= r_data[5530];
                
                r_data[5532] <= r_data[5531];
                
                r_data[5533] <= r_data[5532];
                
                r_data[5534] <= r_data[5533];
                
                r_data[5535] <= r_data[5534];
                
                r_data[5536] <= r_data[5535];
                
                r_data[5537] <= r_data[5536];
                
                r_data[5538] <= r_data[5537];
                
                r_data[5539] <= r_data[5538];
                
                r_data[5540] <= r_data[5539];
                
                r_data[5541] <= r_data[5540];
                
                r_data[5542] <= r_data[5541];
                
                r_data[5543] <= r_data[5542];
                
                r_data[5544] <= r_data[5543];
                
                r_data[5545] <= r_data[5544];
                
                r_data[5546] <= r_data[5545];
                
                r_data[5547] <= r_data[5546];
                
                r_data[5548] <= r_data[5547];
                
                r_data[5549] <= r_data[5548];
                
                r_data[5550] <= r_data[5549];
                
                r_data[5551] <= r_data[5550];
                
                r_data[5552] <= r_data[5551];
                
                r_data[5553] <= r_data[5552];
                
                r_data[5554] <= r_data[5553];
                
                r_data[5555] <= r_data[5554];
                
                r_data[5556] <= r_data[5555];
                
                r_data[5557] <= r_data[5556];
                
                r_data[5558] <= r_data[5557];
                
                r_data[5559] <= r_data[5558];
                
                r_data[5560] <= r_data[5559];
                
                r_data[5561] <= r_data[5560];
                
                r_data[5562] <= r_data[5561];
                
                r_data[5563] <= r_data[5562];
                
                r_data[5564] <= r_data[5563];
                
                r_data[5565] <= r_data[5564];
                
                r_data[5566] <= r_data[5565];
                
                r_data[5567] <= r_data[5566];
                
                r_data[5568] <= r_data[5567];
                
                r_data[5569] <= r_data[5568];
                
                r_data[5570] <= r_data[5569];
                
                r_data[5571] <= r_data[5570];
                
                r_data[5572] <= r_data[5571];
                
                r_data[5573] <= r_data[5572];
                
                r_data[5574] <= r_data[5573];
                
                r_data[5575] <= r_data[5574];
                
                r_data[5576] <= r_data[5575];
                
                r_data[5577] <= r_data[5576];
                
                r_data[5578] <= r_data[5577];
                
                r_data[5579] <= r_data[5578];
                
                r_data[5580] <= r_data[5579];
                
                r_data[5581] <= r_data[5580];
                
                r_data[5582] <= r_data[5581];
                
                r_data[5583] <= r_data[5582];
                
                r_data[5584] <= r_data[5583];
                
                r_data[5585] <= r_data[5584];
                
                r_data[5586] <= r_data[5585];
                
                r_data[5587] <= r_data[5586];
                
                r_data[5588] <= r_data[5587];
                
                r_data[5589] <= r_data[5588];
                
                r_data[5590] <= r_data[5589];
                
                r_data[5591] <= r_data[5590];
                
                r_data[5592] <= r_data[5591];
                
                r_data[5593] <= r_data[5592];
                
                r_data[5594] <= r_data[5593];
                
                r_data[5595] <= r_data[5594];
                
                r_data[5596] <= r_data[5595];
                
                r_data[5597] <= r_data[5596];
                
                r_data[5598] <= r_data[5597];
                
                r_data[5599] <= r_data[5598];
                
                r_data[5600] <= r_data[5599];
                
                r_data[5601] <= r_data[5600];
                
                r_data[5602] <= r_data[5601];
                
                r_data[5603] <= r_data[5602];
                
                r_data[5604] <= r_data[5603];
                
                r_data[5605] <= r_data[5604];
                
                r_data[5606] <= r_data[5605];
                
                r_data[5607] <= r_data[5606];
                
                r_data[5608] <= r_data[5607];
                
                r_data[5609] <= r_data[5608];
                
                r_data[5610] <= r_data[5609];
                
                r_data[5611] <= r_data[5610];
                
                r_data[5612] <= r_data[5611];
                
                r_data[5613] <= r_data[5612];
                
                r_data[5614] <= r_data[5613];
                
                r_data[5615] <= r_data[5614];
                
                r_data[5616] <= r_data[5615];
                
                r_data[5617] <= r_data[5616];
                
                r_data[5618] <= r_data[5617];
                
                r_data[5619] <= r_data[5618];
                
                r_data[5620] <= r_data[5619];
                
                r_data[5621] <= r_data[5620];
                
                r_data[5622] <= r_data[5621];
                
                r_data[5623] <= r_data[5622];
                
                r_data[5624] <= r_data[5623];
                
                r_data[5625] <= r_data[5624];
                
                r_data[5626] <= r_data[5625];
                
                r_data[5627] <= r_data[5626];
                
                r_data[5628] <= r_data[5627];
                
                r_data[5629] <= r_data[5628];
                
                r_data[5630] <= r_data[5629];
                
                r_data[5631] <= r_data[5630];
                
                r_data[5632] <= r_data[5631];
                
                r_data[5633] <= r_data[5632];
                
                r_data[5634] <= r_data[5633];
                
                r_data[5635] <= r_data[5634];
                
                r_data[5636] <= r_data[5635];
                
                r_data[5637] <= r_data[5636];
                
                r_data[5638] <= r_data[5637];
                
                r_data[5639] <= r_data[5638];
                
                r_data[5640] <= r_data[5639];
                
                r_data[5641] <= r_data[5640];
                
                r_data[5642] <= r_data[5641];
                
                r_data[5643] <= r_data[5642];
                
                r_data[5644] <= r_data[5643];
                
                r_data[5645] <= r_data[5644];
                
                r_data[5646] <= r_data[5645];
                
                r_data[5647] <= r_data[5646];
                
                r_data[5648] <= r_data[5647];
                
                r_data[5649] <= r_data[5648];
                
                r_data[5650] <= r_data[5649];
                
                r_data[5651] <= r_data[5650];
                
                r_data[5652] <= r_data[5651];
                
                r_data[5653] <= r_data[5652];
                
                r_data[5654] <= r_data[5653];
                
                r_data[5655] <= r_data[5654];
                
                r_data[5656] <= r_data[5655];
                
                r_data[5657] <= r_data[5656];
                
                r_data[5658] <= r_data[5657];
                
                r_data[5659] <= r_data[5658];
                
                r_data[5660] <= r_data[5659];
                
                r_data[5661] <= r_data[5660];
                
                r_data[5662] <= r_data[5661];
                
                r_data[5663] <= r_data[5662];
                
                r_data[5664] <= r_data[5663];
                
                r_data[5665] <= r_data[5664];
                
                r_data[5666] <= r_data[5665];
                
                r_data[5667] <= r_data[5666];
                
                r_data[5668] <= r_data[5667];
                
                r_data[5669] <= r_data[5668];
                
                r_data[5670] <= r_data[5669];
                
                r_data[5671] <= r_data[5670];
                
                r_data[5672] <= r_data[5671];
                
                r_data[5673] <= r_data[5672];
                
                r_data[5674] <= r_data[5673];
                
                r_data[5675] <= r_data[5674];
                
                r_data[5676] <= r_data[5675];
                
                r_data[5677] <= r_data[5676];
                
                r_data[5678] <= r_data[5677];
                
                r_data[5679] <= r_data[5678];
                
                r_data[5680] <= r_data[5679];
                
                r_data[5681] <= r_data[5680];
                
                r_data[5682] <= r_data[5681];
                
                r_data[5683] <= r_data[5682];
                
                r_data[5684] <= r_data[5683];
                
                r_data[5685] <= r_data[5684];
                
                r_data[5686] <= r_data[5685];
                
                r_data[5687] <= r_data[5686];
                
                r_data[5688] <= r_data[5687];
                
                r_data[5689] <= r_data[5688];
                
                r_data[5690] <= r_data[5689];
                
                r_data[5691] <= r_data[5690];
                
                r_data[5692] <= r_data[5691];
                
                r_data[5693] <= r_data[5692];
                
                r_data[5694] <= r_data[5693];
                
                r_data[5695] <= r_data[5694];
                
                r_data[5696] <= r_data[5695];
                
                r_data[5697] <= r_data[5696];
                
                r_data[5698] <= r_data[5697];
                
                r_data[5699] <= r_data[5698];
                
                r_data[5700] <= r_data[5699];
                
                r_data[5701] <= r_data[5700];
                
                r_data[5702] <= r_data[5701];
                
                r_data[5703] <= r_data[5702];
                
                r_data[5704] <= r_data[5703];
                
                r_data[5705] <= r_data[5704];
                
                r_data[5706] <= r_data[5705];
                
                r_data[5707] <= r_data[5706];
                
                r_data[5708] <= r_data[5707];
                
                r_data[5709] <= r_data[5708];
                
                r_data[5710] <= r_data[5709];
                
                r_data[5711] <= r_data[5710];
                
                r_data[5712] <= r_data[5711];
                
                r_data[5713] <= r_data[5712];
                
                r_data[5714] <= r_data[5713];
                
                r_data[5715] <= r_data[5714];
                
                r_data[5716] <= r_data[5715];
                
                r_data[5717] <= r_data[5716];
                
                r_data[5718] <= r_data[5717];
                
                r_data[5719] <= r_data[5718];
                
                r_data[5720] <= r_data[5719];
                
                r_data[5721] <= r_data[5720];
                
                r_data[5722] <= r_data[5721];
                
                r_data[5723] <= r_data[5722];
                
                r_data[5724] <= r_data[5723];
                
                r_data[5725] <= r_data[5724];
                
                r_data[5726] <= r_data[5725];
                
                r_data[5727] <= r_data[5726];
                
                r_data[5728] <= r_data[5727];
                
                r_data[5729] <= r_data[5728];
                
                r_data[5730] <= r_data[5729];
                
                r_data[5731] <= r_data[5730];
                
                r_data[5732] <= r_data[5731];
                
                r_data[5733] <= r_data[5732];
                
                r_data[5734] <= r_data[5733];
                
                r_data[5735] <= r_data[5734];
                
                r_data[5736] <= r_data[5735];
                
                r_data[5737] <= r_data[5736];
                
                r_data[5738] <= r_data[5737];
                
                r_data[5739] <= r_data[5738];
                
                r_data[5740] <= r_data[5739];
                
                r_data[5741] <= r_data[5740];
                
                r_data[5742] <= r_data[5741];
                
                r_data[5743] <= r_data[5742];
                
                r_data[5744] <= r_data[5743];
                
                r_data[5745] <= r_data[5744];
                
                r_data[5746] <= r_data[5745];
                
                r_data[5747] <= r_data[5746];
                
                r_data[5748] <= r_data[5747];
                
                r_data[5749] <= r_data[5748];
                
                r_data[5750] <= r_data[5749];
                
                r_data[5751] <= r_data[5750];
                
                r_data[5752] <= r_data[5751];
                
                r_data[5753] <= r_data[5752];
                
                r_data[5754] <= r_data[5753];
                
                r_data[5755] <= r_data[5754];
                
                r_data[5756] <= r_data[5755];
                
                r_data[5757] <= r_data[5756];
                
                r_data[5758] <= r_data[5757];
                
                r_data[5759] <= r_data[5758];
                
                r_data[5760] <= r_data[5759];
                
                r_data[5761] <= r_data[5760];
                
                r_data[5762] <= r_data[5761];
                
                r_data[5763] <= r_data[5762];
                
                r_data[5764] <= r_data[5763];
                
                r_data[5765] <= r_data[5764];
                
                r_data[5766] <= r_data[5765];
                
                r_data[5767] <= r_data[5766];
                
                r_data[5768] <= r_data[5767];
                
                r_data[5769] <= r_data[5768];
                
                r_data[5770] <= r_data[5769];
                
                r_data[5771] <= r_data[5770];
                
                r_data[5772] <= r_data[5771];
                
                r_data[5773] <= r_data[5772];
                
                r_data[5774] <= r_data[5773];
                
                r_data[5775] <= r_data[5774];
                
                r_data[5776] <= r_data[5775];
                
                r_data[5777] <= r_data[5776];
                
                r_data[5778] <= r_data[5777];
                
                r_data[5779] <= r_data[5778];
                
                r_data[5780] <= r_data[5779];
                
                r_data[5781] <= r_data[5780];
                
                r_data[5782] <= r_data[5781];
                
                r_data[5783] <= r_data[5782];
                
                r_data[5784] <= r_data[5783];
                
                r_data[5785] <= r_data[5784];
                
                r_data[5786] <= r_data[5785];
                
                r_data[5787] <= r_data[5786];
                
                r_data[5788] <= r_data[5787];
                
                r_data[5789] <= r_data[5788];
                
                r_data[5790] <= r_data[5789];
                
                r_data[5791] <= r_data[5790];
                
                r_data[5792] <= r_data[5791];
                
                r_data[5793] <= r_data[5792];
                
                r_data[5794] <= r_data[5793];
                
                r_data[5795] <= r_data[5794];
                
                r_data[5796] <= r_data[5795];
                
                r_data[5797] <= r_data[5796];
                
                r_data[5798] <= r_data[5797];
                
                r_data[5799] <= r_data[5798];
                
                r_data[5800] <= r_data[5799];
                
                r_data[5801] <= r_data[5800];
                
                r_data[5802] <= r_data[5801];
                
                r_data[5803] <= r_data[5802];
                
                r_data[5804] <= r_data[5803];
                
                r_data[5805] <= r_data[5804];
                
                r_data[5806] <= r_data[5805];
                
                r_data[5807] <= r_data[5806];
                
                r_data[5808] <= r_data[5807];
                
                r_data[5809] <= r_data[5808];
                
                r_data[5810] <= r_data[5809];
                
                r_data[5811] <= r_data[5810];
                
                r_data[5812] <= r_data[5811];
                
                r_data[5813] <= r_data[5812];
                
                r_data[5814] <= r_data[5813];
                
                r_data[5815] <= r_data[5814];
                
                r_data[5816] <= r_data[5815];
                
                r_data[5817] <= r_data[5816];
                
                r_data[5818] <= r_data[5817];
                
                r_data[5819] <= r_data[5818];
                
                r_data[5820] <= r_data[5819];
                
                r_data[5821] <= r_data[5820];
                
                r_data[5822] <= r_data[5821];
                
                r_data[5823] <= r_data[5822];
                
                r_data[5824] <= r_data[5823];
                
                r_data[5825] <= r_data[5824];
                
                r_data[5826] <= r_data[5825];
                
                r_data[5827] <= r_data[5826];
                
                r_data[5828] <= r_data[5827];
                
                r_data[5829] <= r_data[5828];
                
                r_data[5830] <= r_data[5829];
                
                r_data[5831] <= r_data[5830];
                
                r_data[5832] <= r_data[5831];
                
                r_data[5833] <= r_data[5832];
                
                r_data[5834] <= r_data[5833];
                
                r_data[5835] <= r_data[5834];
                
                r_data[5836] <= r_data[5835];
                
                r_data[5837] <= r_data[5836];
                
                r_data[5838] <= r_data[5837];
                
                r_data[5839] <= r_data[5838];
                
                r_data[5840] <= r_data[5839];
                
                r_data[5841] <= r_data[5840];
                
                r_data[5842] <= r_data[5841];
                
                r_data[5843] <= r_data[5842];
                
                r_data[5844] <= r_data[5843];
                
                r_data[5845] <= r_data[5844];
                
                r_data[5846] <= r_data[5845];
                
                r_data[5847] <= r_data[5846];
                
                r_data[5848] <= r_data[5847];
                
                r_data[5849] <= r_data[5848];
                
                r_data[5850] <= r_data[5849];
                
                r_data[5851] <= r_data[5850];
                
                r_data[5852] <= r_data[5851];
                
                r_data[5853] <= r_data[5852];
                
                r_data[5854] <= r_data[5853];
                
                r_data[5855] <= r_data[5854];
                
                r_data[5856] <= r_data[5855];
                
                r_data[5857] <= r_data[5856];
                
                r_data[5858] <= r_data[5857];
                
                r_data[5859] <= r_data[5858];
                
                r_data[5860] <= r_data[5859];
                
                r_data[5861] <= r_data[5860];
                
                r_data[5862] <= r_data[5861];
                
                r_data[5863] <= r_data[5862];
                
                r_data[5864] <= r_data[5863];
                
                r_data[5865] <= r_data[5864];
                
                r_data[5866] <= r_data[5865];
                
                r_data[5867] <= r_data[5866];
                
                r_data[5868] <= r_data[5867];
                
                r_data[5869] <= r_data[5868];
                
                r_data[5870] <= r_data[5869];
                
                r_data[5871] <= r_data[5870];
                
                r_data[5872] <= r_data[5871];
                
                r_data[5873] <= r_data[5872];
                
                r_data[5874] <= r_data[5873];
                
                r_data[5875] <= r_data[5874];
                
                r_data[5876] <= r_data[5875];
                
                r_data[5877] <= r_data[5876];
                
                r_data[5878] <= r_data[5877];
                
                r_data[5879] <= r_data[5878];
                
                r_data[5880] <= r_data[5879];
                
                r_data[5881] <= r_data[5880];
                
                r_data[5882] <= r_data[5881];
                
                r_data[5883] <= r_data[5882];
                
                r_data[5884] <= r_data[5883];
                
                r_data[5885] <= r_data[5884];
                
                r_data[5886] <= r_data[5885];
                
                r_data[5887] <= r_data[5886];
                
                r_data[5888] <= r_data[5887];
                
                r_data[5889] <= r_data[5888];
                
                r_data[5890] <= r_data[5889];
                
                r_data[5891] <= r_data[5890];
                
                r_data[5892] <= r_data[5891];
                
                r_data[5893] <= r_data[5892];
                
                r_data[5894] <= r_data[5893];
                
                r_data[5895] <= r_data[5894];
                
                r_data[5896] <= r_data[5895];
                
                r_data[5897] <= r_data[5896];
                
                r_data[5898] <= r_data[5897];
                
                r_data[5899] <= r_data[5898];
                
                r_data[5900] <= r_data[5899];
                
                r_data[5901] <= r_data[5900];
                
                r_data[5902] <= r_data[5901];
                
                r_data[5903] <= r_data[5902];
                
                r_data[5904] <= r_data[5903];
                
                r_data[5905] <= r_data[5904];
                
                r_data[5906] <= r_data[5905];
                
                r_data[5907] <= r_data[5906];
                
                r_data[5908] <= r_data[5907];
                
                r_data[5909] <= r_data[5908];
                
                r_data[5910] <= r_data[5909];
                
                r_data[5911] <= r_data[5910];
                
                r_data[5912] <= r_data[5911];
                
                r_data[5913] <= r_data[5912];
                
                r_data[5914] <= r_data[5913];
                
                r_data[5915] <= r_data[5914];
                
                r_data[5916] <= r_data[5915];
                
                r_data[5917] <= r_data[5916];
                
                r_data[5918] <= r_data[5917];
                
                r_data[5919] <= r_data[5918];
                
                r_data[5920] <= r_data[5919];
                
                r_data[5921] <= r_data[5920];
                
                r_data[5922] <= r_data[5921];
                
                r_data[5923] <= r_data[5922];
                
                r_data[5924] <= r_data[5923];
                
                r_data[5925] <= r_data[5924];
                
                r_data[5926] <= r_data[5925];
                
                r_data[5927] <= r_data[5926];
                
                r_data[5928] <= r_data[5927];
                
                r_data[5929] <= r_data[5928];
                
                r_data[5930] <= r_data[5929];
                
                r_data[5931] <= r_data[5930];
                
                r_data[5932] <= r_data[5931];
                
                r_data[5933] <= r_data[5932];
                
                r_data[5934] <= r_data[5933];
                
                r_data[5935] <= r_data[5934];
                
                r_data[5936] <= r_data[5935];
                
                r_data[5937] <= r_data[5936];
                
                r_data[5938] <= r_data[5937];
                
                r_data[5939] <= r_data[5938];
                
                r_data[5940] <= r_data[5939];
                
                r_data[5941] <= r_data[5940];
                
                r_data[5942] <= r_data[5941];
                
                r_data[5943] <= r_data[5942];
                
                r_data[5944] <= r_data[5943];
                
                r_data[5945] <= r_data[5944];
                
                r_data[5946] <= r_data[5945];
                
                r_data[5947] <= r_data[5946];
                
                r_data[5948] <= r_data[5947];
                
                r_data[5949] <= r_data[5948];
                
                r_data[5950] <= r_data[5949];
                
                r_data[5951] <= r_data[5950];
                
                r_data[5952] <= r_data[5951];
                
                r_data[5953] <= r_data[5952];
                
                r_data[5954] <= r_data[5953];
                
                r_data[5955] <= r_data[5954];
                
                r_data[5956] <= r_data[5955];
                
                r_data[5957] <= r_data[5956];
                
                r_data[5958] <= r_data[5957];
                
                r_data[5959] <= r_data[5958];
                
                r_data[5960] <= r_data[5959];
                
                r_data[5961] <= r_data[5960];
                
                r_data[5962] <= r_data[5961];
                
                r_data[5963] <= r_data[5962];
                
                r_data[5964] <= r_data[5963];
                
                r_data[5965] <= r_data[5964];
                
                r_data[5966] <= r_data[5965];
                
                r_data[5967] <= r_data[5966];
                
                r_data[5968] <= r_data[5967];
                
                r_data[5969] <= r_data[5968];
                
                r_data[5970] <= r_data[5969];
                
                r_data[5971] <= r_data[5970];
                
                r_data[5972] <= r_data[5971];
                
                r_data[5973] <= r_data[5972];
                
                r_data[5974] <= r_data[5973];
                
                r_data[5975] <= r_data[5974];
                
                r_data[5976] <= r_data[5975];
                
                r_data[5977] <= r_data[5976];
                
                r_data[5978] <= r_data[5977];
                
                r_data[5979] <= r_data[5978];
                
                r_data[5980] <= r_data[5979];
                
                r_data[5981] <= r_data[5980];
                
                r_data[5982] <= r_data[5981];
                
                r_data[5983] <= r_data[5982];
                
                r_data[5984] <= r_data[5983];
                
                r_data[5985] <= r_data[5984];
                
                r_data[5986] <= r_data[5985];
                
                r_data[5987] <= r_data[5986];
                
                r_data[5988] <= r_data[5987];
                
                r_data[5989] <= r_data[5988];
                
                r_data[5990] <= r_data[5989];
                
                r_data[5991] <= r_data[5990];
                
                r_data[5992] <= r_data[5991];
                
                r_data[5993] <= r_data[5992];
                
                r_data[5994] <= r_data[5993];
                
                r_data[5995] <= r_data[5994];
                
                r_data[5996] <= r_data[5995];
                
                r_data[5997] <= r_data[5996];
                
                r_data[5998] <= r_data[5997];
                
                r_data[5999] <= r_data[5998];
                
                r_data[6000] <= r_data[5999];
                
                r_data[6001] <= r_data[6000];
                
                r_data[6002] <= r_data[6001];
                
                r_data[6003] <= r_data[6002];
                
                r_data[6004] <= r_data[6003];
                
                r_data[6005] <= r_data[6004];
                
                r_data[6006] <= r_data[6005];
                
                r_data[6007] <= r_data[6006];
                
                r_data[6008] <= r_data[6007];
                
                r_data[6009] <= r_data[6008];
                
                r_data[6010] <= r_data[6009];
                
                r_data[6011] <= r_data[6010];
                
                r_data[6012] <= r_data[6011];
                
                r_data[6013] <= r_data[6012];
                
                r_data[6014] <= r_data[6013];
                
                r_data[6015] <= r_data[6014];
                
                r_data[6016] <= r_data[6015];
                
                r_data[6017] <= r_data[6016];
                
                r_data[6018] <= r_data[6017];
                
                r_data[6019] <= r_data[6018];
                
                r_data[6020] <= r_data[6019];
                
                r_data[6021] <= r_data[6020];
                
                r_data[6022] <= r_data[6021];
                
                r_data[6023] <= r_data[6022];
                
                r_data[6024] <= r_data[6023];
                
                r_data[6025] <= r_data[6024];
                
                r_data[6026] <= r_data[6025];
                
                r_data[6027] <= r_data[6026];
                
                r_data[6028] <= r_data[6027];
                
                r_data[6029] <= r_data[6028];
                
                r_data[6030] <= r_data[6029];
                
                r_data[6031] <= r_data[6030];
                
                r_data[6032] <= r_data[6031];
                
                r_data[6033] <= r_data[6032];
                
                r_data[6034] <= r_data[6033];
                
                r_data[6035] <= r_data[6034];
                
                r_data[6036] <= r_data[6035];
                
                r_data[6037] <= r_data[6036];
                
                r_data[6038] <= r_data[6037];
                
                r_data[6039] <= r_data[6038];
                
                r_data[6040] <= r_data[6039];
                
                r_data[6041] <= r_data[6040];
                
                r_data[6042] <= r_data[6041];
                
                r_data[6043] <= r_data[6042];
                
                r_data[6044] <= r_data[6043];
                
                r_data[6045] <= r_data[6044];
                
                r_data[6046] <= r_data[6045];
                
                r_data[6047] <= r_data[6046];
                
                r_data[6048] <= r_data[6047];
                
                r_data[6049] <= r_data[6048];
                
                r_data[6050] <= r_data[6049];
                
                r_data[6051] <= r_data[6050];
                
                r_data[6052] <= r_data[6051];
                
                r_data[6053] <= r_data[6052];
                
                r_data[6054] <= r_data[6053];
                
                r_data[6055] <= r_data[6054];
                
                r_data[6056] <= r_data[6055];
                
                r_data[6057] <= r_data[6056];
                
                r_data[6058] <= r_data[6057];
                
                r_data[6059] <= r_data[6058];
                
                r_data[6060] <= r_data[6059];
                
                r_data[6061] <= r_data[6060];
                
                r_data[6062] <= r_data[6061];
                
                r_data[6063] <= r_data[6062];
                
                r_data[6064] <= r_data[6063];
                
                r_data[6065] <= r_data[6064];
                
                r_data[6066] <= r_data[6065];
                
                r_data[6067] <= r_data[6066];
                
                r_data[6068] <= r_data[6067];
                
                r_data[6069] <= r_data[6068];
                
                r_data[6070] <= r_data[6069];
                
                r_data[6071] <= r_data[6070];
                
                r_data[6072] <= r_data[6071];
                
                r_data[6073] <= r_data[6072];
                
                r_data[6074] <= r_data[6073];
                
                r_data[6075] <= r_data[6074];
                
                r_data[6076] <= r_data[6075];
                
                r_data[6077] <= r_data[6076];
                
                r_data[6078] <= r_data[6077];
                
                r_data[6079] <= r_data[6078];
                
                r_data[6080] <= r_data[6079];
                
                r_data[6081] <= r_data[6080];
                
                r_data[6082] <= r_data[6081];
                
                r_data[6083] <= r_data[6082];
                
                r_data[6084] <= r_data[6083];
                
                r_data[6085] <= r_data[6084];
                
                r_data[6086] <= r_data[6085];
                
                r_data[6087] <= r_data[6086];
                
                r_data[6088] <= r_data[6087];
                
                r_data[6089] <= r_data[6088];
                
                r_data[6090] <= r_data[6089];
                
                r_data[6091] <= r_data[6090];
                
                r_data[6092] <= r_data[6091];
                
                r_data[6093] <= r_data[6092];
                
                r_data[6094] <= r_data[6093];
                
                r_data[6095] <= r_data[6094];
                
                r_data[6096] <= r_data[6095];
                
                r_data[6097] <= r_data[6096];
                
                r_data[6098] <= r_data[6097];
                
                r_data[6099] <= r_data[6098];
                
                r_data[6100] <= r_data[6099];
                
                r_data[6101] <= r_data[6100];
                
                r_data[6102] <= r_data[6101];
                
                r_data[6103] <= r_data[6102];
                
                r_data[6104] <= r_data[6103];
                
                r_data[6105] <= r_data[6104];
                
                r_data[6106] <= r_data[6105];
                
                r_data[6107] <= r_data[6106];
                
                r_data[6108] <= r_data[6107];
                
                r_data[6109] <= r_data[6108];
                
                r_data[6110] <= r_data[6109];
                
                r_data[6111] <= r_data[6110];
                
                r_data[6112] <= r_data[6111];
                
                r_data[6113] <= r_data[6112];
                
                r_data[6114] <= r_data[6113];
                
                r_data[6115] <= r_data[6114];
                
                r_data[6116] <= r_data[6115];
                
                r_data[6117] <= r_data[6116];
                
                r_data[6118] <= r_data[6117];
                
                r_data[6119] <= r_data[6118];
                
                r_data[6120] <= r_data[6119];
                
                r_data[6121] <= r_data[6120];
                
                r_data[6122] <= r_data[6121];
                
                r_data[6123] <= r_data[6122];
                
                r_data[6124] <= r_data[6123];
                
                r_data[6125] <= r_data[6124];
                
                r_data[6126] <= r_data[6125];
                
                r_data[6127] <= r_data[6126];
                
                r_data[6128] <= r_data[6127];
                
                r_data[6129] <= r_data[6128];
                
                r_data[6130] <= r_data[6129];
                
                r_data[6131] <= r_data[6130];
                
                r_data[6132] <= r_data[6131];
                
                r_data[6133] <= r_data[6132];
                
                r_data[6134] <= r_data[6133];
                
                r_data[6135] <= r_data[6134];
                
                r_data[6136] <= r_data[6135];
                
                r_data[6137] <= r_data[6136];
                
                r_data[6138] <= r_data[6137];
                
                r_data[6139] <= r_data[6138];
                
                r_data[6140] <= r_data[6139];
                
                r_data[6141] <= r_data[6140];
                
                r_data[6142] <= r_data[6141];
                
                r_data[6143] <= r_data[6142];
                
                r_data[6144] <= r_data[6143];
                
                r_data[6145] <= r_data[6144];
                
                r_data[6146] <= r_data[6145];
                
                r_data[6147] <= r_data[6146];
                
                r_data[6148] <= r_data[6147];
                
                r_data[6149] <= r_data[6148];
                
                r_data[6150] <= r_data[6149];
                
                r_data[6151] <= r_data[6150];
                
                r_data[6152] <= r_data[6151];
                
                r_data[6153] <= r_data[6152];
                
                r_data[6154] <= r_data[6153];
                
                r_data[6155] <= r_data[6154];
                
                r_data[6156] <= r_data[6155];
                
                r_data[6157] <= r_data[6156];
                
                r_data[6158] <= r_data[6157];
                
                r_data[6159] <= r_data[6158];
                
                r_data[6160] <= r_data[6159];
                
                r_data[6161] <= r_data[6160];
                
                r_data[6162] <= r_data[6161];
                
                r_data[6163] <= r_data[6162];
                
                r_data[6164] <= r_data[6163];
                
                r_data[6165] <= r_data[6164];
                
                r_data[6166] <= r_data[6165];
                
                r_data[6167] <= r_data[6166];
                
                r_data[6168] <= r_data[6167];
                
                r_data[6169] <= r_data[6168];
                
                r_data[6170] <= r_data[6169];
                
                r_data[6171] <= r_data[6170];
                
                r_data[6172] <= r_data[6171];
                
                r_data[6173] <= r_data[6172];
                
                r_data[6174] <= r_data[6173];
                
                r_data[6175] <= r_data[6174];
                
                r_data[6176] <= r_data[6175];
                
                r_data[6177] <= r_data[6176];
                
                r_data[6178] <= r_data[6177];
                
                r_data[6179] <= r_data[6178];
                
                r_data[6180] <= r_data[6179];
                
                r_data[6181] <= r_data[6180];
                
                r_data[6182] <= r_data[6181];
                
                r_data[6183] <= r_data[6182];
                
                r_data[6184] <= r_data[6183];
                
                r_data[6185] <= r_data[6184];
                
                r_data[6186] <= r_data[6185];
                
                r_data[6187] <= r_data[6186];
                
                r_data[6188] <= r_data[6187];
                
                r_data[6189] <= r_data[6188];
                
                r_data[6190] <= r_data[6189];
                
                r_data[6191] <= r_data[6190];
                
                r_data[6192] <= r_data[6191];
                
                r_data[6193] <= r_data[6192];
                
                r_data[6194] <= r_data[6193];
                
                r_data[6195] <= r_data[6194];
                
                r_data[6196] <= r_data[6195];
                
                r_data[6197] <= r_data[6196];
                
                r_data[6198] <= r_data[6197];
                
                r_data[6199] <= r_data[6198];
                
                r_data[6200] <= r_data[6199];
                
                r_data[6201] <= r_data[6200];
                
                r_data[6202] <= r_data[6201];
                
                r_data[6203] <= r_data[6202];
                
                r_data[6204] <= r_data[6203];
                
                r_data[6205] <= r_data[6204];
                
                r_data[6206] <= r_data[6205];
                
                r_data[6207] <= r_data[6206];
                
                r_data[6208] <= r_data[6207];
                
                r_data[6209] <= r_data[6208];
                
                r_data[6210] <= r_data[6209];
                
                r_data[6211] <= r_data[6210];
                
                r_data[6212] <= r_data[6211];
                
                r_data[6213] <= r_data[6212];
                
                r_data[6214] <= r_data[6213];
                
                r_data[6215] <= r_data[6214];
                
                r_data[6216] <= r_data[6215];
                
                r_data[6217] <= r_data[6216];
                
                r_data[6218] <= r_data[6217];
                
                r_data[6219] <= r_data[6218];
                
                r_data[6220] <= r_data[6219];
                
                r_data[6221] <= r_data[6220];
                
                r_data[6222] <= r_data[6221];
                
                r_data[6223] <= r_data[6222];
                
                r_data[6224] <= r_data[6223];
                
                r_data[6225] <= r_data[6224];
                
                r_data[6226] <= r_data[6225];
                
                r_data[6227] <= r_data[6226];
                
                r_data[6228] <= r_data[6227];
                
                r_data[6229] <= r_data[6228];
                
                r_data[6230] <= r_data[6229];
                
                r_data[6231] <= r_data[6230];
                
                r_data[6232] <= r_data[6231];
                
                r_data[6233] <= r_data[6232];
                
                r_data[6234] <= r_data[6233];
                
                r_data[6235] <= r_data[6234];
                
                r_data[6236] <= r_data[6235];
                
                r_data[6237] <= r_data[6236];
                
                r_data[6238] <= r_data[6237];
                
                r_data[6239] <= r_data[6238];
                
                r_data[6240] <= r_data[6239];
                
                r_data[6241] <= r_data[6240];
                
                r_data[6242] <= r_data[6241];
                
                r_data[6243] <= r_data[6242];
                
                r_data[6244] <= r_data[6243];
                
                r_data[6245] <= r_data[6244];
                
                r_data[6246] <= r_data[6245];
                
                r_data[6247] <= r_data[6246];
                
                r_data[6248] <= r_data[6247];
                
                r_data[6249] <= r_data[6248];
                
                r_data[6250] <= r_data[6249];
                
                r_data[6251] <= r_data[6250];
                
                r_data[6252] <= r_data[6251];
                
                r_data[6253] <= r_data[6252];
                
                r_data[6254] <= r_data[6253];
                
                r_data[6255] <= r_data[6254];
                
                r_data[6256] <= r_data[6255];
                
                r_data[6257] <= r_data[6256];
                
                r_data[6258] <= r_data[6257];
                
                r_data[6259] <= r_data[6258];
                
                r_data[6260] <= r_data[6259];
                
                r_data[6261] <= r_data[6260];
                
                r_data[6262] <= r_data[6261];
                
                r_data[6263] <= r_data[6262];
                
                r_data[6264] <= r_data[6263];
                
                r_data[6265] <= r_data[6264];
                
                r_data[6266] <= r_data[6265];
                
                r_data[6267] <= r_data[6266];
                
                r_data[6268] <= r_data[6267];
                
                r_data[6269] <= r_data[6268];
                
                r_data[6270] <= r_data[6269];
                
                r_data[6271] <= r_data[6270];
                
                r_data[6272] <= r_data[6271];
                
                r_data[6273] <= r_data[6272];
                
                r_data[6274] <= r_data[6273];
                
                r_data[6275] <= r_data[6274];
                
                r_data[6276] <= r_data[6275];
                
                r_data[6277] <= r_data[6276];
                
                r_data[6278] <= r_data[6277];
                
                r_data[6279] <= r_data[6278];
                
                r_data[6280] <= r_data[6279];
                
                r_data[6281] <= r_data[6280];
                
                r_data[6282] <= r_data[6281];
                
                r_data[6283] <= r_data[6282];
                
                r_data[6284] <= r_data[6283];
                
                r_data[6285] <= r_data[6284];
                
                r_data[6286] <= r_data[6285];
                
                r_data[6287] <= r_data[6286];
                
                r_data[6288] <= r_data[6287];
                
                r_data[6289] <= r_data[6288];
                
                r_data[6290] <= r_data[6289];
                
                r_data[6291] <= r_data[6290];
                
                r_data[6292] <= r_data[6291];
                
                r_data[6293] <= r_data[6292];
                
                r_data[6294] <= r_data[6293];
                
                r_data[6295] <= r_data[6294];
                
                r_data[6296] <= r_data[6295];
                
                r_data[6297] <= r_data[6296];
                
                r_data[6298] <= r_data[6297];
                
                r_data[6299] <= r_data[6298];
                
                r_data[6300] <= r_data[6299];
                
                r_data[6301] <= r_data[6300];
                
                r_data[6302] <= r_data[6301];
                
                r_data[6303] <= r_data[6302];
                
                r_data[6304] <= r_data[6303];
                
                r_data[6305] <= r_data[6304];
                
                r_data[6306] <= r_data[6305];
                
                r_data[6307] <= r_data[6306];
                
                r_data[6308] <= r_data[6307];
                
                r_data[6309] <= r_data[6308];
                
                r_data[6310] <= r_data[6309];
                
                r_data[6311] <= r_data[6310];
                
                r_data[6312] <= r_data[6311];
                
                r_data[6313] <= r_data[6312];
                
                r_data[6314] <= r_data[6313];
                
                r_data[6315] <= r_data[6314];
                
                r_data[6316] <= r_data[6315];
                
                r_data[6317] <= r_data[6316];
                
                r_data[6318] <= r_data[6317];
                
                r_data[6319] <= r_data[6318];
                
                r_data[6320] <= r_data[6319];
                
                r_data[6321] <= r_data[6320];
                
                r_data[6322] <= r_data[6321];
                
                r_data[6323] <= r_data[6322];
                
                r_data[6324] <= r_data[6323];
                
                r_data[6325] <= r_data[6324];
                
                r_data[6326] <= r_data[6325];
                
                r_data[6327] <= r_data[6326];
                
                r_data[6328] <= r_data[6327];
                
                r_data[6329] <= r_data[6328];
                
                r_data[6330] <= r_data[6329];
                
                r_data[6331] <= r_data[6330];
                
                r_data[6332] <= r_data[6331];
                
                r_data[6333] <= r_data[6332];
                
                r_data[6334] <= r_data[6333];
                
                r_data[6335] <= r_data[6334];
                
                r_data[6336] <= r_data[6335];
                
                r_data[6337] <= r_data[6336];
                
                r_data[6338] <= r_data[6337];
                
                r_data[6339] <= r_data[6338];
                
                r_data[6340] <= r_data[6339];
                
                r_data[6341] <= r_data[6340];
                
                r_data[6342] <= r_data[6341];
                
                r_data[6343] <= r_data[6342];
                
                r_data[6344] <= r_data[6343];
                
                r_data[6345] <= r_data[6344];
                
                r_data[6346] <= r_data[6345];
                
                r_data[6347] <= r_data[6346];
                
                r_data[6348] <= r_data[6347];
                
                r_data[6349] <= r_data[6348];
                
                r_data[6350] <= r_data[6349];
                
                r_data[6351] <= r_data[6350];
                
                r_data[6352] <= r_data[6351];
                
                r_data[6353] <= r_data[6352];
                
                r_data[6354] <= r_data[6353];
                
                r_data[6355] <= r_data[6354];
                
                r_data[6356] <= r_data[6355];
                
                r_data[6357] <= r_data[6356];
                
                r_data[6358] <= r_data[6357];
                
                r_data[6359] <= r_data[6358];
                
                r_data[6360] <= r_data[6359];
                
                r_data[6361] <= r_data[6360];
                
                r_data[6362] <= r_data[6361];
                
                r_data[6363] <= r_data[6362];
                
                r_data[6364] <= r_data[6363];
                
                r_data[6365] <= r_data[6364];
                
                r_data[6366] <= r_data[6365];
                
                r_data[6367] <= r_data[6366];
                
                r_data[6368] <= r_data[6367];
                
                r_data[6369] <= r_data[6368];
                
                r_data[6370] <= r_data[6369];
                
                r_data[6371] <= r_data[6370];
                
                r_data[6372] <= r_data[6371];
                
                r_data[6373] <= r_data[6372];
                
                r_data[6374] <= r_data[6373];
                
                r_data[6375] <= r_data[6374];
                
                r_data[6376] <= r_data[6375];
                
                r_data[6377] <= r_data[6376];
                
                r_data[6378] <= r_data[6377];
                
                r_data[6379] <= r_data[6378];
                
                r_data[6380] <= r_data[6379];
                
                r_data[6381] <= r_data[6380];
                
                r_data[6382] <= r_data[6381];
                
                r_data[6383] <= r_data[6382];
                
                r_data[6384] <= r_data[6383];
                
                r_data[6385] <= r_data[6384];
                
                r_data[6386] <= r_data[6385];
                
                r_data[6387] <= r_data[6386];
                
                r_data[6388] <= r_data[6387];
                
                r_data[6389] <= r_data[6388];
                
                r_data[6390] <= r_data[6389];
                
                r_data[6391] <= r_data[6390];
                
                r_data[6392] <= r_data[6391];
                
                r_data[6393] <= r_data[6392];
                
                r_data[6394] <= r_data[6393];
                
                r_data[6395] <= r_data[6394];
                
                r_data[6396] <= r_data[6395];
                
                r_data[6397] <= r_data[6396];
                
                r_data[6398] <= r_data[6397];
                
                r_data[6399] <= r_data[6398];
                
                r_data[6400] <= r_data[6399];
                
                r_data[6401] <= r_data[6400];
                
                r_data[6402] <= r_data[6401];
                
                r_data[6403] <= r_data[6402];
                
                r_data[6404] <= r_data[6403];
                
                r_data[6405] <= r_data[6404];
                
                r_data[6406] <= r_data[6405];
                
                r_data[6407] <= r_data[6406];
                
                r_data[6408] <= r_data[6407];
                
                r_data[6409] <= r_data[6408];
                
                r_data[6410] <= r_data[6409];
                
                r_data[6411] <= r_data[6410];
                
                r_data[6412] <= r_data[6411];
                
                r_data[6413] <= r_data[6412];
                
                r_data[6414] <= r_data[6413];
                
                r_data[6415] <= r_data[6414];
                
                r_data[6416] <= r_data[6415];
                
                r_data[6417] <= r_data[6416];
                
                r_data[6418] <= r_data[6417];
                
                r_data[6419] <= r_data[6418];
                
                r_data[6420] <= r_data[6419];
                
                r_data[6421] <= r_data[6420];
                
                r_data[6422] <= r_data[6421];
                
                r_data[6423] <= r_data[6422];
                
                r_data[6424] <= r_data[6423];
                
                r_data[6425] <= r_data[6424];
                
                r_data[6426] <= r_data[6425];
                
                r_data[6427] <= r_data[6426];
                
                r_data[6428] <= r_data[6427];
                
                r_data[6429] <= r_data[6428];
                
                r_data[6430] <= r_data[6429];
                
                r_data[6431] <= r_data[6430];
                
                r_data[6432] <= r_data[6431];
                
                r_data[6433] <= r_data[6432];
                
                r_data[6434] <= r_data[6433];
                
                r_data[6435] <= r_data[6434];
                
                r_data[6436] <= r_data[6435];
                
                r_data[6437] <= r_data[6436];
                
                r_data[6438] <= r_data[6437];
                
                r_data[6439] <= r_data[6438];
                
                r_data[6440] <= r_data[6439];
                
                r_data[6441] <= r_data[6440];
                
                r_data[6442] <= r_data[6441];
                
                r_data[6443] <= r_data[6442];
                
                r_data[6444] <= r_data[6443];
                
                r_data[6445] <= r_data[6444];
                
                r_data[6446] <= r_data[6445];
                
                r_data[6447] <= r_data[6446];
                
                r_data[6448] <= r_data[6447];
                
                r_data[6449] <= r_data[6448];
                
                r_data[6450] <= r_data[6449];
                
                r_data[6451] <= r_data[6450];
                
                r_data[6452] <= r_data[6451];
                
                r_data[6453] <= r_data[6452];
                
                r_data[6454] <= r_data[6453];
                
                r_data[6455] <= r_data[6454];
                
                r_data[6456] <= r_data[6455];
                
                r_data[6457] <= r_data[6456];
                
                r_data[6458] <= r_data[6457];
                
                r_data[6459] <= r_data[6458];
                
                r_data[6460] <= r_data[6459];
                
                r_data[6461] <= r_data[6460];
                
                r_data[6462] <= r_data[6461];
                
                r_data[6463] <= r_data[6462];
                
                r_data[6464] <= r_data[6463];
                
                r_data[6465] <= r_data[6464];
                
                r_data[6466] <= r_data[6465];
                
                r_data[6467] <= r_data[6466];
                
                r_data[6468] <= r_data[6467];
                
                r_data[6469] <= r_data[6468];
                
                r_data[6470] <= r_data[6469];
                
                r_data[6471] <= r_data[6470];
                
                r_data[6472] <= r_data[6471];
                
                r_data[6473] <= r_data[6472];
                
                r_data[6474] <= r_data[6473];
                
                r_data[6475] <= r_data[6474];
                
                r_data[6476] <= r_data[6475];
                
                r_data[6477] <= r_data[6476];
                
                r_data[6478] <= r_data[6477];
                
                r_data[6479] <= r_data[6478];
                
                r_data[6480] <= r_data[6479];
                
                r_data[6481] <= r_data[6480];
                
                r_data[6482] <= r_data[6481];
                
                r_data[6483] <= r_data[6482];
                
                r_data[6484] <= r_data[6483];
                
                r_data[6485] <= r_data[6484];
                
                r_data[6486] <= r_data[6485];
                
                r_data[6487] <= r_data[6486];
                
                r_data[6488] <= r_data[6487];
                
                r_data[6489] <= r_data[6488];
                
                r_data[6490] <= r_data[6489];
                
                r_data[6491] <= r_data[6490];
                
                r_data[6492] <= r_data[6491];
                
                r_data[6493] <= r_data[6492];
                
                r_data[6494] <= r_data[6493];
                
                r_data[6495] <= r_data[6494];
                
                r_data[6496] <= r_data[6495];
                
                r_data[6497] <= r_data[6496];
                
                r_data[6498] <= r_data[6497];
                
                r_data[6499] <= r_data[6498];
                
                r_data[6500] <= r_data[6499];
                
                r_data[6501] <= r_data[6500];
                
                r_data[6502] <= r_data[6501];
                
                r_data[6503] <= r_data[6502];
                
                r_data[6504] <= r_data[6503];
                
                r_data[6505] <= r_data[6504];
                
                r_data[6506] <= r_data[6505];
                
                r_data[6507] <= r_data[6506];
                
                r_data[6508] <= r_data[6507];
                
                r_data[6509] <= r_data[6508];
                
                r_data[6510] <= r_data[6509];
                
                r_data[6511] <= r_data[6510];
                
                r_data[6512] <= r_data[6511];
                
                r_data[6513] <= r_data[6512];
                
                r_data[6514] <= r_data[6513];
                
                r_data[6515] <= r_data[6514];
                
                r_data[6516] <= r_data[6515];
                
                r_data[6517] <= r_data[6516];
                
                r_data[6518] <= r_data[6517];
                
                r_data[6519] <= r_data[6518];
                
                r_data[6520] <= r_data[6519];
                
                r_data[6521] <= r_data[6520];
                
                r_data[6522] <= r_data[6521];
                
                r_data[6523] <= r_data[6522];
                
                r_data[6524] <= r_data[6523];
                
                r_data[6525] <= r_data[6524];
                
                r_data[6526] <= r_data[6525];
                
                r_data[6527] <= r_data[6526];
                
                r_data[6528] <= r_data[6527];
                
                r_data[6529] <= r_data[6528];
                
                r_data[6530] <= r_data[6529];
                
                r_data[6531] <= r_data[6530];
                
                r_data[6532] <= r_data[6531];
                
                r_data[6533] <= r_data[6532];
                
                r_data[6534] <= r_data[6533];
                
                r_data[6535] <= r_data[6534];
                
                r_data[6536] <= r_data[6535];
                
                r_data[6537] <= r_data[6536];
                
                r_data[6538] <= r_data[6537];
                
                r_data[6539] <= r_data[6538];
                
                r_data[6540] <= r_data[6539];
                
                r_data[6541] <= r_data[6540];
                
                r_data[6542] <= r_data[6541];
                
                r_data[6543] <= r_data[6542];
                
                r_data[6544] <= r_data[6543];
                
                r_data[6545] <= r_data[6544];
                
                r_data[6546] <= r_data[6545];
                
                r_data[6547] <= r_data[6546];
                
                r_data[6548] <= r_data[6547];
                
                r_data[6549] <= r_data[6548];
                
                r_data[6550] <= r_data[6549];
                
                r_data[6551] <= r_data[6550];
                
                r_data[6552] <= r_data[6551];
                
                r_data[6553] <= r_data[6552];
                
                r_data[6554] <= r_data[6553];
                
                r_data[6555] <= r_data[6554];
                
                r_data[6556] <= r_data[6555];
                
                r_data[6557] <= r_data[6556];
                
                r_data[6558] <= r_data[6557];
                
                r_data[6559] <= r_data[6558];
                
                r_data[6560] <= r_data[6559];
                
                r_data[6561] <= r_data[6560];
                
                r_data[6562] <= r_data[6561];
                
                r_data[6563] <= r_data[6562];
                
                r_data[6564] <= r_data[6563];
                
                r_data[6565] <= r_data[6564];
                
                r_data[6566] <= r_data[6565];
                
                r_data[6567] <= r_data[6566];
                
                r_data[6568] <= r_data[6567];
                
                r_data[6569] <= r_data[6568];
                
                r_data[6570] <= r_data[6569];
                
                r_data[6571] <= r_data[6570];
                
                r_data[6572] <= r_data[6571];
                
                r_data[6573] <= r_data[6572];
                
                r_data[6574] <= r_data[6573];
                
                r_data[6575] <= r_data[6574];
                
                r_data[6576] <= r_data[6575];
                
                r_data[6577] <= r_data[6576];
                
                r_data[6578] <= r_data[6577];
                
                r_data[6579] <= r_data[6578];
                
                r_data[6580] <= r_data[6579];
                
                r_data[6581] <= r_data[6580];
                
                r_data[6582] <= r_data[6581];
                
                r_data[6583] <= r_data[6582];
                
                r_data[6584] <= r_data[6583];
                
                r_data[6585] <= r_data[6584];
                
                r_data[6586] <= r_data[6585];
                
                r_data[6587] <= r_data[6586];
                
                r_data[6588] <= r_data[6587];
                
                r_data[6589] <= r_data[6588];
                
                r_data[6590] <= r_data[6589];
                
                r_data[6591] <= r_data[6590];
                
                r_data[6592] <= r_data[6591];
                
                r_data[6593] <= r_data[6592];
                
                r_data[6594] <= r_data[6593];
                
                r_data[6595] <= r_data[6594];
                
                r_data[6596] <= r_data[6595];
                
                r_data[6597] <= r_data[6596];
                
                r_data[6598] <= r_data[6597];
                
                r_data[6599] <= r_data[6598];
                
                r_data[6600] <= r_data[6599];
                
                r_data[6601] <= r_data[6600];
                
                r_data[6602] <= r_data[6601];
                
                r_data[6603] <= r_data[6602];
                
                r_data[6604] <= r_data[6603];
                
                r_data[6605] <= r_data[6604];
                
                r_data[6606] <= r_data[6605];
                
                r_data[6607] <= r_data[6606];
                
                r_data[6608] <= r_data[6607];
                
                r_data[6609] <= r_data[6608];
                
                r_data[6610] <= r_data[6609];
                
                r_data[6611] <= r_data[6610];
                
                r_data[6612] <= r_data[6611];
                
                r_data[6613] <= r_data[6612];
                
                r_data[6614] <= r_data[6613];
                
                r_data[6615] <= r_data[6614];
                
                r_data[6616] <= r_data[6615];
                
                r_data[6617] <= r_data[6616];
                
                r_data[6618] <= r_data[6617];
                
                r_data[6619] <= r_data[6618];
                
                r_data[6620] <= r_data[6619];
                
                r_data[6621] <= r_data[6620];
                
                r_data[6622] <= r_data[6621];
                
                r_data[6623] <= r_data[6622];
                
                r_data[6624] <= r_data[6623];
                
                r_data[6625] <= r_data[6624];
                
                r_data[6626] <= r_data[6625];
                
                r_data[6627] <= r_data[6626];
                
                r_data[6628] <= r_data[6627];
                
                r_data[6629] <= r_data[6628];
                
                r_data[6630] <= r_data[6629];
                
                r_data[6631] <= r_data[6630];
                
                r_data[6632] <= r_data[6631];
                
                r_data[6633] <= r_data[6632];
                
                r_data[6634] <= r_data[6633];
                
                r_data[6635] <= r_data[6634];
                
                r_data[6636] <= r_data[6635];
                
                r_data[6637] <= r_data[6636];
                
                r_data[6638] <= r_data[6637];
                
                r_data[6639] <= r_data[6638];
                
                r_data[6640] <= r_data[6639];
                
                r_data[6641] <= r_data[6640];
                
                r_data[6642] <= r_data[6641];
                
                r_data[6643] <= r_data[6642];
                
                r_data[6644] <= r_data[6643];
                
                r_data[6645] <= r_data[6644];
                
                r_data[6646] <= r_data[6645];
                
                r_data[6647] <= r_data[6646];
                
                r_data[6648] <= r_data[6647];
                
                r_data[6649] <= r_data[6648];
                
                r_data[6650] <= r_data[6649];
                
                r_data[6651] <= r_data[6650];
                
                r_data[6652] <= r_data[6651];
                
                r_data[6653] <= r_data[6652];
                
                r_data[6654] <= r_data[6653];
                
                r_data[6655] <= r_data[6654];
                
                r_data[6656] <= r_data[6655];
                
                r_data[6657] <= r_data[6656];
                
                r_data[6658] <= r_data[6657];
                
                r_data[6659] <= r_data[6658];
                
                r_data[6660] <= r_data[6659];
                
                r_data[6661] <= r_data[6660];
                
                r_data[6662] <= r_data[6661];
                
                r_data[6663] <= r_data[6662];
                
                r_data[6664] <= r_data[6663];
                
                r_data[6665] <= r_data[6664];
                
                r_data[6666] <= r_data[6665];
                
                r_data[6667] <= r_data[6666];
                
                r_data[6668] <= r_data[6667];
                
                r_data[6669] <= r_data[6668];
                
                r_data[6670] <= r_data[6669];
                
                r_data[6671] <= r_data[6670];
                
                r_data[6672] <= r_data[6671];
                
                r_data[6673] <= r_data[6672];
                
                r_data[6674] <= r_data[6673];
                
                r_data[6675] <= r_data[6674];
                
                r_data[6676] <= r_data[6675];
                
                r_data[6677] <= r_data[6676];
                
                r_data[6678] <= r_data[6677];
                
                r_data[6679] <= r_data[6678];
                
                r_data[6680] <= r_data[6679];
                
                r_data[6681] <= r_data[6680];
                
                r_data[6682] <= r_data[6681];
                
                r_data[6683] <= r_data[6682];
                
                r_data[6684] <= r_data[6683];
                
                r_data[6685] <= r_data[6684];
                
                r_data[6686] <= r_data[6685];
                
                r_data[6687] <= r_data[6686];
                
                r_data[6688] <= r_data[6687];
                
                r_data[6689] <= r_data[6688];
                
                r_data[6690] <= r_data[6689];
                
                r_data[6691] <= r_data[6690];
                
                r_data[6692] <= r_data[6691];
                
                r_data[6693] <= r_data[6692];
                
                r_data[6694] <= r_data[6693];
                
                r_data[6695] <= r_data[6694];
                
                r_data[6696] <= r_data[6695];
                
                r_data[6697] <= r_data[6696];
                
                r_data[6698] <= r_data[6697];
                
                r_data[6699] <= r_data[6698];
                
                r_data[6700] <= r_data[6699];
                
                r_data[6701] <= r_data[6700];
                
                r_data[6702] <= r_data[6701];
                
                r_data[6703] <= r_data[6702];
                
                r_data[6704] <= r_data[6703];
                
                r_data[6705] <= r_data[6704];
                
                r_data[6706] <= r_data[6705];
                
                r_data[6707] <= r_data[6706];
                
                r_data[6708] <= r_data[6707];
                
                r_data[6709] <= r_data[6708];
                
                r_data[6710] <= r_data[6709];
                
                r_data[6711] <= r_data[6710];
                
                r_data[6712] <= r_data[6711];
                
                r_data[6713] <= r_data[6712];
                
                r_data[6714] <= r_data[6713];
                
                r_data[6715] <= r_data[6714];
                
                r_data[6716] <= r_data[6715];
                
                r_data[6717] <= r_data[6716];
                
                r_data[6718] <= r_data[6717];
                
                r_data[6719] <= r_data[6718];
                
                r_data[6720] <= r_data[6719];
                
                r_data[6721] <= r_data[6720];
                
                r_data[6722] <= r_data[6721];
                
                r_data[6723] <= r_data[6722];
                
                r_data[6724] <= r_data[6723];
                
                r_data[6725] <= r_data[6724];
                
                r_data[6726] <= r_data[6725];
                
                r_data[6727] <= r_data[6726];
                
                r_data[6728] <= r_data[6727];
                
                r_data[6729] <= r_data[6728];
                
                r_data[6730] <= r_data[6729];
                
                r_data[6731] <= r_data[6730];
                
                r_data[6732] <= r_data[6731];
                
                r_data[6733] <= r_data[6732];
                
                r_data[6734] <= r_data[6733];
                
                r_data[6735] <= r_data[6734];
                
                r_data[6736] <= r_data[6735];
                
                r_data[6737] <= r_data[6736];
                
                r_data[6738] <= r_data[6737];
                
                r_data[6739] <= r_data[6738];
                
                r_data[6740] <= r_data[6739];
                
                r_data[6741] <= r_data[6740];
                
                r_data[6742] <= r_data[6741];
                
                r_data[6743] <= r_data[6742];
                
                r_data[6744] <= r_data[6743];
                
                r_data[6745] <= r_data[6744];
                
                r_data[6746] <= r_data[6745];
                
                r_data[6747] <= r_data[6746];
                
                r_data[6748] <= r_data[6747];
                
                r_data[6749] <= r_data[6748];
                
                r_data[6750] <= r_data[6749];
                
                r_data[6751] <= r_data[6750];
                
                r_data[6752] <= r_data[6751];
                
                r_data[6753] <= r_data[6752];
                
                r_data[6754] <= r_data[6753];
                
                r_data[6755] <= r_data[6754];
                
                r_data[6756] <= r_data[6755];
                
                r_data[6757] <= r_data[6756];
                
                r_data[6758] <= r_data[6757];
                
                r_data[6759] <= r_data[6758];
                
                r_data[6760] <= r_data[6759];
                
                r_data[6761] <= r_data[6760];
                
                r_data[6762] <= r_data[6761];
                
                r_data[6763] <= r_data[6762];
                
                r_data[6764] <= r_data[6763];
                
                r_data[6765] <= r_data[6764];
                
                r_data[6766] <= r_data[6765];
                
                r_data[6767] <= r_data[6766];
                
                r_data[6768] <= r_data[6767];
                
                r_data[6769] <= r_data[6768];
                
                r_data[6770] <= r_data[6769];
                
                r_data[6771] <= r_data[6770];
                
                r_data[6772] <= r_data[6771];
                
                r_data[6773] <= r_data[6772];
                
                r_data[6774] <= r_data[6773];
                
                r_data[6775] <= r_data[6774];
                
                r_data[6776] <= r_data[6775];
                
                r_data[6777] <= r_data[6776];
                
                r_data[6778] <= r_data[6777];
                
                r_data[6779] <= r_data[6778];
                
                r_data[6780] <= r_data[6779];
                
                r_data[6781] <= r_data[6780];
                
                r_data[6782] <= r_data[6781];
                
                r_data[6783] <= r_data[6782];
                
                r_data[6784] <= r_data[6783];
                
                r_data[6785] <= r_data[6784];
                
                r_data[6786] <= r_data[6785];
                
                r_data[6787] <= r_data[6786];
                
                r_data[6788] <= r_data[6787];
                
                r_data[6789] <= r_data[6788];
                
                r_data[6790] <= r_data[6789];
                
                r_data[6791] <= r_data[6790];
                
                r_data[6792] <= r_data[6791];
                
                r_data[6793] <= r_data[6792];
                
                r_data[6794] <= r_data[6793];
                
                r_data[6795] <= r_data[6794];
                
                r_data[6796] <= r_data[6795];
                
                r_data[6797] <= r_data[6796];
                
                r_data[6798] <= r_data[6797];
                
                r_data[6799] <= r_data[6798];
                
                r_data[6800] <= r_data[6799];
                
                r_data[6801] <= r_data[6800];
                
                r_data[6802] <= r_data[6801];
                
                r_data[6803] <= r_data[6802];
                
                r_data[6804] <= r_data[6803];
                
                r_data[6805] <= r_data[6804];
                
                r_data[6806] <= r_data[6805];
                
                r_data[6807] <= r_data[6806];
                
                r_data[6808] <= r_data[6807];
                
                r_data[6809] <= r_data[6808];
                
                r_data[6810] <= r_data[6809];
                
                r_data[6811] <= r_data[6810];
                
                r_data[6812] <= r_data[6811];
                
                r_data[6813] <= r_data[6812];
                
                r_data[6814] <= r_data[6813];
                
                r_data[6815] <= r_data[6814];
                
                r_data[6816] <= r_data[6815];
                
                r_data[6817] <= r_data[6816];
                
                r_data[6818] <= r_data[6817];
                
                r_data[6819] <= r_data[6818];
                
                r_data[6820] <= r_data[6819];
                
                r_data[6821] <= r_data[6820];
                
                r_data[6822] <= r_data[6821];
                
                r_data[6823] <= r_data[6822];
                
                r_data[6824] <= r_data[6823];
                
                r_data[6825] <= r_data[6824];
                
                r_data[6826] <= r_data[6825];
                
                r_data[6827] <= r_data[6826];
                
                r_data[6828] <= r_data[6827];
                
                r_data[6829] <= r_data[6828];
                
                r_data[6830] <= r_data[6829];
                
                r_data[6831] <= r_data[6830];
                
                r_data[6832] <= r_data[6831];
                
                r_data[6833] <= r_data[6832];
                
                r_data[6834] <= r_data[6833];
                
                r_data[6835] <= r_data[6834];
                
                r_data[6836] <= r_data[6835];
                
                r_data[6837] <= r_data[6836];
                
                r_data[6838] <= r_data[6837];
                
                r_data[6839] <= r_data[6838];
                
                r_data[6840] <= r_data[6839];
                
                r_data[6841] <= r_data[6840];
                
                r_data[6842] <= r_data[6841];
                
                r_data[6843] <= r_data[6842];
                
                r_data[6844] <= r_data[6843];
                
                r_data[6845] <= r_data[6844];
                
                r_data[6846] <= r_data[6845];
                
                r_data[6847] <= r_data[6846];
                
                r_data[6848] <= r_data[6847];
                
                r_data[6849] <= r_data[6848];
                
                r_data[6850] <= r_data[6849];
                
                r_data[6851] <= r_data[6850];
                
                r_data[6852] <= r_data[6851];
                
                r_data[6853] <= r_data[6852];
                
                r_data[6854] <= r_data[6853];
                
                r_data[6855] <= r_data[6854];
                
                r_data[6856] <= r_data[6855];
                
                r_data[6857] <= r_data[6856];
                
                r_data[6858] <= r_data[6857];
                
                r_data[6859] <= r_data[6858];
                
                r_data[6860] <= r_data[6859];
                
                r_data[6861] <= r_data[6860];
                
                r_data[6862] <= r_data[6861];
                
                r_data[6863] <= r_data[6862];
                
                r_data[6864] <= r_data[6863];
                
                r_data[6865] <= r_data[6864];
                
                r_data[6866] <= r_data[6865];
                
                r_data[6867] <= r_data[6866];
                
                r_data[6868] <= r_data[6867];
                
                r_data[6869] <= r_data[6868];
                
                r_data[6870] <= r_data[6869];
                
                r_data[6871] <= r_data[6870];
                
                r_data[6872] <= r_data[6871];
                
                r_data[6873] <= r_data[6872];
                
                r_data[6874] <= r_data[6873];
                
                r_data[6875] <= r_data[6874];
                
                r_data[6876] <= r_data[6875];
                
                r_data[6877] <= r_data[6876];
                
                r_data[6878] <= r_data[6877];
                
                r_data[6879] <= r_data[6878];
                
                r_data[6880] <= r_data[6879];
                
                r_data[6881] <= r_data[6880];
                
                r_data[6882] <= r_data[6881];
                
                r_data[6883] <= r_data[6882];
                
                r_data[6884] <= r_data[6883];
                
                r_data[6885] <= r_data[6884];
                
                r_data[6886] <= r_data[6885];
                
                r_data[6887] <= r_data[6886];
                
                r_data[6888] <= r_data[6887];
                
                r_data[6889] <= r_data[6888];
                
                r_data[6890] <= r_data[6889];
                
                r_data[6891] <= r_data[6890];
                
                r_data[6892] <= r_data[6891];
                
                r_data[6893] <= r_data[6892];
                
                r_data[6894] <= r_data[6893];
                
                r_data[6895] <= r_data[6894];
                
                r_data[6896] <= r_data[6895];
                
                r_data[6897] <= r_data[6896];
                
                r_data[6898] <= r_data[6897];
                
                r_data[6899] <= r_data[6898];
                
                r_data[6900] <= r_data[6899];
                
                r_data[6901] <= r_data[6900];
                
                r_data[6902] <= r_data[6901];
                
                r_data[6903] <= r_data[6902];
                
                r_data[6904] <= r_data[6903];
                
                r_data[6905] <= r_data[6904];
                
                r_data[6906] <= r_data[6905];
                
                r_data[6907] <= r_data[6906];
                
                r_data[6908] <= r_data[6907];
                
                r_data[6909] <= r_data[6908];
                
                r_data[6910] <= r_data[6909];
                
                r_data[6911] <= r_data[6910];
                
                r_data[6912] <= r_data[6911];
                
                r_data[6913] <= r_data[6912];
                
                r_data[6914] <= r_data[6913];
                
                r_data[6915] <= r_data[6914];
                
                r_data[6916] <= r_data[6915];
                
                r_data[6917] <= r_data[6916];
                
                r_data[6918] <= r_data[6917];
                
                r_data[6919] <= r_data[6918];
                
                r_data[6920] <= r_data[6919];
                
                r_data[6921] <= r_data[6920];
                
                r_data[6922] <= r_data[6921];
                
                r_data[6923] <= r_data[6922];
                
                r_data[6924] <= r_data[6923];
                
                r_data[6925] <= r_data[6924];
                
                r_data[6926] <= r_data[6925];
                
                r_data[6927] <= r_data[6926];
                
                r_data[6928] <= r_data[6927];
                
                r_data[6929] <= r_data[6928];
                
                r_data[6930] <= r_data[6929];
                
                r_data[6931] <= r_data[6930];
                
                r_data[6932] <= r_data[6931];
                
                r_data[6933] <= r_data[6932];
                
                r_data[6934] <= r_data[6933];
                
                r_data[6935] <= r_data[6934];
                
                r_data[6936] <= r_data[6935];
                
                r_data[6937] <= r_data[6936];
                
                r_data[6938] <= r_data[6937];
                
                r_data[6939] <= r_data[6938];
                
                r_data[6940] <= r_data[6939];
                
                r_data[6941] <= r_data[6940];
                
                r_data[6942] <= r_data[6941];
                
                r_data[6943] <= r_data[6942];
                
                r_data[6944] <= r_data[6943];
                
                r_data[6945] <= r_data[6944];
                
                r_data[6946] <= r_data[6945];
                
                r_data[6947] <= r_data[6946];
                
                r_data[6948] <= r_data[6947];
                
                r_data[6949] <= r_data[6948];
                
                r_data[6950] <= r_data[6949];
                
                r_data[6951] <= r_data[6950];
                
                r_data[6952] <= r_data[6951];
                
                r_data[6953] <= r_data[6952];
                
                r_data[6954] <= r_data[6953];
                
                r_data[6955] <= r_data[6954];
                
                r_data[6956] <= r_data[6955];
                
                r_data[6957] <= r_data[6956];
                
                r_data[6958] <= r_data[6957];
                
                r_data[6959] <= r_data[6958];
                
                r_data[6960] <= r_data[6959];
                
                r_data[6961] <= r_data[6960];
                
                r_data[6962] <= r_data[6961];
                
                r_data[6963] <= r_data[6962];
                
                r_data[6964] <= r_data[6963];
                
                r_data[6965] <= r_data[6964];
                
                r_data[6966] <= r_data[6965];
                
                r_data[6967] <= r_data[6966];
                
                r_data[6968] <= r_data[6967];
                
                r_data[6969] <= r_data[6968];
                
                r_data[6970] <= r_data[6969];
                
                r_data[6971] <= r_data[6970];
                
                r_data[6972] <= r_data[6971];
                
                r_data[6973] <= r_data[6972];
                
                r_data[6974] <= r_data[6973];
                
                r_data[6975] <= r_data[6974];
                
                r_data[6976] <= r_data[6975];
                
                r_data[6977] <= r_data[6976];
                
                r_data[6978] <= r_data[6977];
                
                r_data[6979] <= r_data[6978];
                
                r_data[6980] <= r_data[6979];
                
                r_data[6981] <= r_data[6980];
                
                r_data[6982] <= r_data[6981];
                
                r_data[6983] <= r_data[6982];
                
                r_data[6984] <= r_data[6983];
                
                r_data[6985] <= r_data[6984];
                
                r_data[6986] <= r_data[6985];
                
                r_data[6987] <= r_data[6986];
                
                r_data[6988] <= r_data[6987];
                
                r_data[6989] <= r_data[6988];
                
                r_data[6990] <= r_data[6989];
                
                r_data[6991] <= r_data[6990];
                
                r_data[6992] <= r_data[6991];
                
                r_data[6993] <= r_data[6992];
                
                r_data[6994] <= r_data[6993];
                
                r_data[6995] <= r_data[6994];
                
                r_data[6996] <= r_data[6995];
                
                r_data[6997] <= r_data[6996];
                
                r_data[6998] <= r_data[6997];
                
                r_data[6999] <= r_data[6998];
                
                r_data[7000] <= r_data[6999];
                
                r_data[7001] <= r_data[7000];
                
                r_data[7002] <= r_data[7001];
                
                r_data[7003] <= r_data[7002];
                
                r_data[7004] <= r_data[7003];
                
                r_data[7005] <= r_data[7004];
                
                r_data[7006] <= r_data[7005];
                
                r_data[7007] <= r_data[7006];
                
                r_data[7008] <= r_data[7007];
                
                r_data[7009] <= r_data[7008];
                
                r_data[7010] <= r_data[7009];
                
                r_data[7011] <= r_data[7010];
                
                r_data[7012] <= r_data[7011];
                
                r_data[7013] <= r_data[7012];
                
                r_data[7014] <= r_data[7013];
                
                r_data[7015] <= r_data[7014];
                
                r_data[7016] <= r_data[7015];
                
                r_data[7017] <= r_data[7016];
                
                r_data[7018] <= r_data[7017];
                
                r_data[7019] <= r_data[7018];
                
                r_data[7020] <= r_data[7019];
                
                r_data[7021] <= r_data[7020];
                
                r_data[7022] <= r_data[7021];
                
                r_data[7023] <= r_data[7022];
                
                r_data[7024] <= r_data[7023];
                
                r_data[7025] <= r_data[7024];
                
                r_data[7026] <= r_data[7025];
                
                r_data[7027] <= r_data[7026];
                
                r_data[7028] <= r_data[7027];
                
                r_data[7029] <= r_data[7028];
                
                r_data[7030] <= r_data[7029];
                
                r_data[7031] <= r_data[7030];
                
                r_data[7032] <= r_data[7031];
                
                r_data[7033] <= r_data[7032];
                
                r_data[7034] <= r_data[7033];
                
                r_data[7035] <= r_data[7034];
                
                r_data[7036] <= r_data[7035];
                
                r_data[7037] <= r_data[7036];
                
                r_data[7038] <= r_data[7037];
                
                r_data[7039] <= r_data[7038];
                
                r_data[7040] <= r_data[7039];
                
                r_data[7041] <= r_data[7040];
                
                r_data[7042] <= r_data[7041];
                
                r_data[7043] <= r_data[7042];
                
                r_data[7044] <= r_data[7043];
                
                r_data[7045] <= r_data[7044];
                
                r_data[7046] <= r_data[7045];
                
                r_data[7047] <= r_data[7046];
                
                r_data[7048] <= r_data[7047];
                
                r_data[7049] <= r_data[7048];
                
                r_data[7050] <= r_data[7049];
                
                r_data[7051] <= r_data[7050];
                
                r_data[7052] <= r_data[7051];
                
                r_data[7053] <= r_data[7052];
                
                r_data[7054] <= r_data[7053];
                
                r_data[7055] <= r_data[7054];
                
                r_data[7056] <= r_data[7055];
                
                r_data[7057] <= r_data[7056];
                
                r_data[7058] <= r_data[7057];
                
                r_data[7059] <= r_data[7058];
                
                r_data[7060] <= r_data[7059];
                
                r_data[7061] <= r_data[7060];
                
                r_data[7062] <= r_data[7061];
                
                r_data[7063] <= r_data[7062];
                
                r_data[7064] <= r_data[7063];
                
                r_data[7065] <= r_data[7064];
                
                r_data[7066] <= r_data[7065];
                
                r_data[7067] <= r_data[7066];
                
                r_data[7068] <= r_data[7067];
                
                r_data[7069] <= r_data[7068];
                
                r_data[7070] <= r_data[7069];
                
                r_data[7071] <= r_data[7070];
                
                r_data[7072] <= r_data[7071];
                
                r_data[7073] <= r_data[7072];
                
                r_data[7074] <= r_data[7073];
                
                r_data[7075] <= r_data[7074];
                
                r_data[7076] <= r_data[7075];
                
                r_data[7077] <= r_data[7076];
                
                r_data[7078] <= r_data[7077];
                
                r_data[7079] <= r_data[7078];
                
                r_data[7080] <= r_data[7079];
                
                r_data[7081] <= r_data[7080];
                
                r_data[7082] <= r_data[7081];
                
                r_data[7083] <= r_data[7082];
                
                r_data[7084] <= r_data[7083];
                
                r_data[7085] <= r_data[7084];
                
                r_data[7086] <= r_data[7085];
                
                r_data[7087] <= r_data[7086];
                
                r_data[7088] <= r_data[7087];
                
                r_data[7089] <= r_data[7088];
                
                r_data[7090] <= r_data[7089];
                
                r_data[7091] <= r_data[7090];
                
                r_data[7092] <= r_data[7091];
                
                r_data[7093] <= r_data[7092];
                
                r_data[7094] <= r_data[7093];
                
                r_data[7095] <= r_data[7094];
                
                r_data[7096] <= r_data[7095];
                
                r_data[7097] <= r_data[7096];
                
                r_data[7098] <= r_data[7097];
                
                r_data[7099] <= r_data[7098];
                
                r_data[7100] <= r_data[7099];
                
                r_data[7101] <= r_data[7100];
                
                r_data[7102] <= r_data[7101];
                
                r_data[7103] <= r_data[7102];
                
                r_data[7104] <= r_data[7103];
                
                r_data[7105] <= r_data[7104];
                
                r_data[7106] <= r_data[7105];
                
                r_data[7107] <= r_data[7106];
                
                r_data[7108] <= r_data[7107];
                
                r_data[7109] <= r_data[7108];
                
                r_data[7110] <= r_data[7109];
                
                r_data[7111] <= r_data[7110];
                
                r_data[7112] <= r_data[7111];
                
                r_data[7113] <= r_data[7112];
                
                r_data[7114] <= r_data[7113];
                
                r_data[7115] <= r_data[7114];
                
                r_data[7116] <= r_data[7115];
                
                r_data[7117] <= r_data[7116];
                
                r_data[7118] <= r_data[7117];
                
                r_data[7119] <= r_data[7118];
                
                r_data[7120] <= r_data[7119];
                
                r_data[7121] <= r_data[7120];
                
                r_data[7122] <= r_data[7121];
                
                r_data[7123] <= r_data[7122];
                
                r_data[7124] <= r_data[7123];
                
                r_data[7125] <= r_data[7124];
                
                r_data[7126] <= r_data[7125];
                
                r_data[7127] <= r_data[7126];
                
                r_data[7128] <= r_data[7127];
                
                r_data[7129] <= r_data[7128];
                
                r_data[7130] <= r_data[7129];
                
                r_data[7131] <= r_data[7130];
                
                r_data[7132] <= r_data[7131];
                
                r_data[7133] <= r_data[7132];
                
                r_data[7134] <= r_data[7133];
                
                r_data[7135] <= r_data[7134];
                
                r_data[7136] <= r_data[7135];
                
                r_data[7137] <= r_data[7136];
                
                r_data[7138] <= r_data[7137];
                
                r_data[7139] <= r_data[7138];
                
                r_data[7140] <= r_data[7139];
                
                r_data[7141] <= r_data[7140];
                
                r_data[7142] <= r_data[7141];
                
                r_data[7143] <= r_data[7142];
                
                r_data[7144] <= r_data[7143];
                
                r_data[7145] <= r_data[7144];
                
                r_data[7146] <= r_data[7145];
                
                r_data[7147] <= r_data[7146];
                
                r_data[7148] <= r_data[7147];
                
                r_data[7149] <= r_data[7148];
                
                r_data[7150] <= r_data[7149];
                
                r_data[7151] <= r_data[7150];
                
                r_data[7152] <= r_data[7151];
                
                r_data[7153] <= r_data[7152];
                
                r_data[7154] <= r_data[7153];
                
                r_data[7155] <= r_data[7154];
                
                r_data[7156] <= r_data[7155];
                
                r_data[7157] <= r_data[7156];
                
                r_data[7158] <= r_data[7157];
                
                r_data[7159] <= r_data[7158];
                
                r_data[7160] <= r_data[7159];
                
                r_data[7161] <= r_data[7160];
                
                r_data[7162] <= r_data[7161];
                
                r_data[7163] <= r_data[7162];
                
                r_data[7164] <= r_data[7163];
                
                r_data[7165] <= r_data[7164];
                
                r_data[7166] <= r_data[7165];
                
                r_data[7167] <= r_data[7166];
                
                r_data[7168] <= r_data[7167];
                
                r_data[7169] <= r_data[7168];
                
                r_data[7170] <= r_data[7169];
                
                r_data[7171] <= r_data[7170];
                
                r_data[7172] <= r_data[7171];
                
                r_data[7173] <= r_data[7172];
                
                r_data[7174] <= r_data[7173];
                
                r_data[7175] <= r_data[7174];
                
                r_data[7176] <= r_data[7175];
                
                r_data[7177] <= r_data[7176];
                
                r_data[7178] <= r_data[7177];
                
                r_data[7179] <= r_data[7178];
                
                r_data[7180] <= r_data[7179];
                
                r_data[7181] <= r_data[7180];
                
                r_data[7182] <= r_data[7181];
                
                r_data[7183] <= r_data[7182];
                
                r_data[7184] <= r_data[7183];
                
                r_data[7185] <= r_data[7184];
                
                r_data[7186] <= r_data[7185];
                
                r_data[7187] <= r_data[7186];
                
                r_data[7188] <= r_data[7187];
                
                r_data[7189] <= r_data[7188];
                
                r_data[7190] <= r_data[7189];
                
                r_data[7191] <= r_data[7190];
                
                r_data[7192] <= r_data[7191];
                
                r_data[7193] <= r_data[7192];
                
                r_data[7194] <= r_data[7193];
                
                r_data[7195] <= r_data[7194];
                
                r_data[7196] <= r_data[7195];
                
                r_data[7197] <= r_data[7196];
                
                r_data[7198] <= r_data[7197];
                
                r_data[7199] <= r_data[7198];
                
                r_data[7200] <= r_data[7199];
                
                r_data[7201] <= r_data[7200];
                
                r_data[7202] <= r_data[7201];
                
                r_data[7203] <= r_data[7202];
                
                r_data[7204] <= r_data[7203];
                
                r_data[7205] <= r_data[7204];
                
                r_data[7206] <= r_data[7205];
                
                r_data[7207] <= r_data[7206];
                
                r_data[7208] <= r_data[7207];
                
                r_data[7209] <= r_data[7208];
                
                r_data[7210] <= r_data[7209];
                
                r_data[7211] <= r_data[7210];
                
                r_data[7212] <= r_data[7211];
                
                r_data[7213] <= r_data[7212];
                
                r_data[7214] <= r_data[7213];
                
                r_data[7215] <= r_data[7214];
                
                r_data[7216] <= r_data[7215];
                
                r_data[7217] <= r_data[7216];
                
                r_data[7218] <= r_data[7217];
                
                r_data[7219] <= r_data[7218];
                
                r_data[7220] <= r_data[7219];
                
                r_data[7221] <= r_data[7220];
                
                r_data[7222] <= r_data[7221];
                
                r_data[7223] <= r_data[7222];
                
                r_data[7224] <= r_data[7223];
                
                r_data[7225] <= r_data[7224];
                
                r_data[7226] <= r_data[7225];
                
                r_data[7227] <= r_data[7226];
                
                r_data[7228] <= r_data[7227];
                
                r_data[7229] <= r_data[7228];
                
                r_data[7230] <= r_data[7229];
                
                r_data[7231] <= r_data[7230];
                
                r_data[7232] <= r_data[7231];
                
                r_data[7233] <= r_data[7232];
                
                r_data[7234] <= r_data[7233];
                
                r_data[7235] <= r_data[7234];
                
                r_data[7236] <= r_data[7235];
                
                r_data[7237] <= r_data[7236];
                
                r_data[7238] <= r_data[7237];
                
                r_data[7239] <= r_data[7238];
                
                r_data[7240] <= r_data[7239];
                
                r_data[7241] <= r_data[7240];
                
                r_data[7242] <= r_data[7241];
                
                r_data[7243] <= r_data[7242];
                
                r_data[7244] <= r_data[7243];
                
                r_data[7245] <= r_data[7244];
                
                r_data[7246] <= r_data[7245];
                
                r_data[7247] <= r_data[7246];
                
                r_data[7248] <= r_data[7247];
                
                r_data[7249] <= r_data[7248];
                
                r_data[7250] <= r_data[7249];
                
                r_data[7251] <= r_data[7250];
                
                r_data[7252] <= r_data[7251];
                
                r_data[7253] <= r_data[7252];
                
                r_data[7254] <= r_data[7253];
                
                r_data[7255] <= r_data[7254];
                
                r_data[7256] <= r_data[7255];
                
                r_data[7257] <= r_data[7256];
                
                r_data[7258] <= r_data[7257];
                
                r_data[7259] <= r_data[7258];
                
                r_data[7260] <= r_data[7259];
                
                r_data[7261] <= r_data[7260];
                
                r_data[7262] <= r_data[7261];
                
                r_data[7263] <= r_data[7262];
                
                r_data[7264] <= r_data[7263];
                
                r_data[7265] <= r_data[7264];
                
                r_data[7266] <= r_data[7265];
                
                r_data[7267] <= r_data[7266];
                
                r_data[7268] <= r_data[7267];
                
                r_data[7269] <= r_data[7268];
                
                r_data[7270] <= r_data[7269];
                
                r_data[7271] <= r_data[7270];
                
                r_data[7272] <= r_data[7271];
                
                r_data[7273] <= r_data[7272];
                
                r_data[7274] <= r_data[7273];
                
                r_data[7275] <= r_data[7274];
                
                r_data[7276] <= r_data[7275];
                
                r_data[7277] <= r_data[7276];
                
                r_data[7278] <= r_data[7277];
                
                r_data[7279] <= r_data[7278];
                
                r_data[7280] <= r_data[7279];
                
                r_data[7281] <= r_data[7280];
                
                r_data[7282] <= r_data[7281];
                
                r_data[7283] <= r_data[7282];
                
                r_data[7284] <= r_data[7283];
                
                r_data[7285] <= r_data[7284];
                
                r_data[7286] <= r_data[7285];
                
                r_data[7287] <= r_data[7286];
                
                r_data[7288] <= r_data[7287];
                
                r_data[7289] <= r_data[7288];
                
                r_data[7290] <= r_data[7289];
                
                r_data[7291] <= r_data[7290];
                
                r_data[7292] <= r_data[7291];
                
                r_data[7293] <= r_data[7292];
                
                r_data[7294] <= r_data[7293];
                
                r_data[7295] <= r_data[7294];
                
                r_data[7296] <= r_data[7295];
                
                r_data[7297] <= r_data[7296];
                
                r_data[7298] <= r_data[7297];
                
                r_data[7299] <= r_data[7298];
                
                r_data[7300] <= r_data[7299];
                
                r_data[7301] <= r_data[7300];
                
                r_data[7302] <= r_data[7301];
                
                r_data[7303] <= r_data[7302];
                
                r_data[7304] <= r_data[7303];
                
                r_data[7305] <= r_data[7304];
                
                r_data[7306] <= r_data[7305];
                
                r_data[7307] <= r_data[7306];
                
                r_data[7308] <= r_data[7307];
                
                r_data[7309] <= r_data[7308];
                
                r_data[7310] <= r_data[7309];
                
                r_data[7311] <= r_data[7310];
                
                r_data[7312] <= r_data[7311];
                
                r_data[7313] <= r_data[7312];
                
                r_data[7314] <= r_data[7313];
                
                r_data[7315] <= r_data[7314];
                
                r_data[7316] <= r_data[7315];
                
                r_data[7317] <= r_data[7316];
                
                r_data[7318] <= r_data[7317];
                
                r_data[7319] <= r_data[7318];
                
                r_data[7320] <= r_data[7319];
                
                r_data[7321] <= r_data[7320];
                
                r_data[7322] <= r_data[7321];
                
                r_data[7323] <= r_data[7322];
                
                r_data[7324] <= r_data[7323];
                
                r_data[7325] <= r_data[7324];
                
                r_data[7326] <= r_data[7325];
                
                r_data[7327] <= r_data[7326];
                
                r_data[7328] <= r_data[7327];
                
                r_data[7329] <= r_data[7328];
                
                r_data[7330] <= r_data[7329];
                
                r_data[7331] <= r_data[7330];
                
                r_data[7332] <= r_data[7331];
                
                r_data[7333] <= r_data[7332];
                
                r_data[7334] <= r_data[7333];
                
                r_data[7335] <= r_data[7334];
                
                r_data[7336] <= r_data[7335];
                
                r_data[7337] <= r_data[7336];
                
                r_data[7338] <= r_data[7337];
                
                r_data[7339] <= r_data[7338];
                
                r_data[7340] <= r_data[7339];
                
                r_data[7341] <= r_data[7340];
                
                r_data[7342] <= r_data[7341];
                
                r_data[7343] <= r_data[7342];
                
                r_data[7344] <= r_data[7343];
                
                r_data[7345] <= r_data[7344];
                
                r_data[7346] <= r_data[7345];
                
                r_data[7347] <= r_data[7346];
                
                r_data[7348] <= r_data[7347];
                
                r_data[7349] <= r_data[7348];
                
                r_data[7350] <= r_data[7349];
                
                r_data[7351] <= r_data[7350];
                
                r_data[7352] <= r_data[7351];
                
                r_data[7353] <= r_data[7352];
                
                r_data[7354] <= r_data[7353];
                
                r_data[7355] <= r_data[7354];
                
                r_data[7356] <= r_data[7355];
                
                r_data[7357] <= r_data[7356];
                
                r_data[7358] <= r_data[7357];
                
                r_data[7359] <= r_data[7358];
                
                r_data[7360] <= r_data[7359];
                
                r_data[7361] <= r_data[7360];
                
                r_data[7362] <= r_data[7361];
                
                r_data[7363] <= r_data[7362];
                
                r_data[7364] <= r_data[7363];
                
                r_data[7365] <= r_data[7364];
                
                r_data[7366] <= r_data[7365];
                
                r_data[7367] <= r_data[7366];
                
                r_data[7368] <= r_data[7367];
                
                r_data[7369] <= r_data[7368];
                
                r_data[7370] <= r_data[7369];
                
                r_data[7371] <= r_data[7370];
                
                r_data[7372] <= r_data[7371];
                
                r_data[7373] <= r_data[7372];
                
                r_data[7374] <= r_data[7373];
                
                r_data[7375] <= r_data[7374];
                
                r_data[7376] <= r_data[7375];
                
                r_data[7377] <= r_data[7376];
                
                r_data[7378] <= r_data[7377];
                
                r_data[7379] <= r_data[7378];
                
                r_data[7380] <= r_data[7379];
                
                r_data[7381] <= r_data[7380];
                
                r_data[7382] <= r_data[7381];
                
                r_data[7383] <= r_data[7382];
                
                r_data[7384] <= r_data[7383];
                
                r_data[7385] <= r_data[7384];
                
                r_data[7386] <= r_data[7385];
                
                r_data[7387] <= r_data[7386];
                
                r_data[7388] <= r_data[7387];
                
                r_data[7389] <= r_data[7388];
                
                r_data[7390] <= r_data[7389];
                
                r_data[7391] <= r_data[7390];
                
                r_data[7392] <= r_data[7391];
                
                r_data[7393] <= r_data[7392];
                
                r_data[7394] <= r_data[7393];
                
                r_data[7395] <= r_data[7394];
                
                r_data[7396] <= r_data[7395];
                
                r_data[7397] <= r_data[7396];
                
                r_data[7398] <= r_data[7397];
                
                r_data[7399] <= r_data[7398];
                
                r_data[7400] <= r_data[7399];
                
                r_data[7401] <= r_data[7400];
                
                r_data[7402] <= r_data[7401];
                
                r_data[7403] <= r_data[7402];
                
                r_data[7404] <= r_data[7403];
                
                r_data[7405] <= r_data[7404];
                
                r_data[7406] <= r_data[7405];
                
                r_data[7407] <= r_data[7406];
                
                r_data[7408] <= r_data[7407];
                
                r_data[7409] <= r_data[7408];
                
                r_data[7410] <= r_data[7409];
                
                r_data[7411] <= r_data[7410];
                
                r_data[7412] <= r_data[7411];
                
                r_data[7413] <= r_data[7412];
                
                r_data[7414] <= r_data[7413];
                
                r_data[7415] <= r_data[7414];
                
                r_data[7416] <= r_data[7415];
                
                r_data[7417] <= r_data[7416];
                
                r_data[7418] <= r_data[7417];
                
                r_data[7419] <= r_data[7418];
                
                r_data[7420] <= r_data[7419];
                
                r_data[7421] <= r_data[7420];
                
                r_data[7422] <= r_data[7421];
                
                r_data[7423] <= r_data[7422];
                
                r_data[7424] <= r_data[7423];
                
                r_data[7425] <= r_data[7424];
                
                r_data[7426] <= r_data[7425];
                
                r_data[7427] <= r_data[7426];
                
                r_data[7428] <= r_data[7427];
                
                r_data[7429] <= r_data[7428];
                
                r_data[7430] <= r_data[7429];
                
                r_data[7431] <= r_data[7430];
                
                r_data[7432] <= r_data[7431];
                
                r_data[7433] <= r_data[7432];
                
                r_data[7434] <= r_data[7433];
                
                r_data[7435] <= r_data[7434];
                
                r_data[7436] <= r_data[7435];
                
                r_data[7437] <= r_data[7436];
                
                r_data[7438] <= r_data[7437];
                
                r_data[7439] <= r_data[7438];
                
                r_data[7440] <= r_data[7439];
                
                r_data[7441] <= r_data[7440];
                
                r_data[7442] <= r_data[7441];
                
                r_data[7443] <= r_data[7442];
                
                r_data[7444] <= r_data[7443];
                
                r_data[7445] <= r_data[7444];
                
                r_data[7446] <= r_data[7445];
                
                r_data[7447] <= r_data[7446];
                
                r_data[7448] <= r_data[7447];
                
                r_data[7449] <= r_data[7448];
                
                r_data[7450] <= r_data[7449];
                
                r_data[7451] <= r_data[7450];
                
                r_data[7452] <= r_data[7451];
                
                r_data[7453] <= r_data[7452];
                
                r_data[7454] <= r_data[7453];
                
                r_data[7455] <= r_data[7454];
                
                r_data[7456] <= r_data[7455];
                
                r_data[7457] <= r_data[7456];
                
                r_data[7458] <= r_data[7457];
                
                r_data[7459] <= r_data[7458];
                
                r_data[7460] <= r_data[7459];
                
                r_data[7461] <= r_data[7460];
                
                r_data[7462] <= r_data[7461];
                
                r_data[7463] <= r_data[7462];
                
                r_data[7464] <= r_data[7463];
                
                r_data[7465] <= r_data[7464];
                
                r_data[7466] <= r_data[7465];
                
                r_data[7467] <= r_data[7466];
                
                r_data[7468] <= r_data[7467];
                
                r_data[7469] <= r_data[7468];
                
                r_data[7470] <= r_data[7469];
                
                r_data[7471] <= r_data[7470];
                
                r_data[7472] <= r_data[7471];
                
                r_data[7473] <= r_data[7472];
                
                r_data[7474] <= r_data[7473];
                
                r_data[7475] <= r_data[7474];
                
                r_data[7476] <= r_data[7475];
                
                r_data[7477] <= r_data[7476];
                
                r_data[7478] <= r_data[7477];
                
                r_data[7479] <= r_data[7478];
                
                r_data[7480] <= r_data[7479];
                
                r_data[7481] <= r_data[7480];
                
                r_data[7482] <= r_data[7481];
                
                r_data[7483] <= r_data[7482];
                
                r_data[7484] <= r_data[7483];
                
                r_data[7485] <= r_data[7484];
                
                r_data[7486] <= r_data[7485];
                
                r_data[7487] <= r_data[7486];
                
                r_data[7488] <= r_data[7487];
                
                r_data[7489] <= r_data[7488];
                
                r_data[7490] <= r_data[7489];
                
                r_data[7491] <= r_data[7490];
                
                r_data[7492] <= r_data[7491];
                
                r_data[7493] <= r_data[7492];
                
                r_data[7494] <= r_data[7493];
                
                r_data[7495] <= r_data[7494];
                
                r_data[7496] <= r_data[7495];
                
                r_data[7497] <= r_data[7496];
                
                r_data[7498] <= r_data[7497];
                
                r_data[7499] <= r_data[7498];
                
                r_data[7500] <= r_data[7499];
                
                r_data[7501] <= r_data[7500];
                
                r_data[7502] <= r_data[7501];
                
                r_data[7503] <= r_data[7502];
                
                r_data[7504] <= r_data[7503];
                
                r_data[7505] <= r_data[7504];
                
                r_data[7506] <= r_data[7505];
                
                r_data[7507] <= r_data[7506];
                
                r_data[7508] <= r_data[7507];
                
                r_data[7509] <= r_data[7508];
                
                r_data[7510] <= r_data[7509];
                
                r_data[7511] <= r_data[7510];
                
                r_data[7512] <= r_data[7511];
                
                r_data[7513] <= r_data[7512];
                
                r_data[7514] <= r_data[7513];
                
                r_data[7515] <= r_data[7514];
                
                r_data[7516] <= r_data[7515];
                
                r_data[7517] <= r_data[7516];
                
                r_data[7518] <= r_data[7517];
                
                r_data[7519] <= r_data[7518];
                
                r_data[7520] <= r_data[7519];
                
                r_data[7521] <= r_data[7520];
                
                r_data[7522] <= r_data[7521];
                
                r_data[7523] <= r_data[7522];
                
                r_data[7524] <= r_data[7523];
                
                r_data[7525] <= r_data[7524];
                
                r_data[7526] <= r_data[7525];
                
                r_data[7527] <= r_data[7526];
                
                r_data[7528] <= r_data[7527];
                
                r_data[7529] <= r_data[7528];
                
                r_data[7530] <= r_data[7529];
                
                r_data[7531] <= r_data[7530];
                
                r_data[7532] <= r_data[7531];
                
                r_data[7533] <= r_data[7532];
                
                r_data[7534] <= r_data[7533];
                
                r_data[7535] <= r_data[7534];
                
                r_data[7536] <= r_data[7535];
                
                r_data[7537] <= r_data[7536];
                
                r_data[7538] <= r_data[7537];
                
                r_data[7539] <= r_data[7538];
                
                r_data[7540] <= r_data[7539];
                
                r_data[7541] <= r_data[7540];
                
                r_data[7542] <= r_data[7541];
                
                r_data[7543] <= r_data[7542];
                
                r_data[7544] <= r_data[7543];
                
                r_data[7545] <= r_data[7544];
                
                r_data[7546] <= r_data[7545];
                
                r_data[7547] <= r_data[7546];
                
                r_data[7548] <= r_data[7547];
                
                r_data[7549] <= r_data[7548];
                
                r_data[7550] <= r_data[7549];
                
                r_data[7551] <= r_data[7550];
                
                r_data[7552] <= r_data[7551];
                
                r_data[7553] <= r_data[7552];
                
                r_data[7554] <= r_data[7553];
                
                r_data[7555] <= r_data[7554];
                
                r_data[7556] <= r_data[7555];
                
                r_data[7557] <= r_data[7556];
                
                r_data[7558] <= r_data[7557];
                
                r_data[7559] <= r_data[7558];
                
                r_data[7560] <= r_data[7559];
                
                r_data[7561] <= r_data[7560];
                
                r_data[7562] <= r_data[7561];
                
                r_data[7563] <= r_data[7562];
                
                r_data[7564] <= r_data[7563];
                
                r_data[7565] <= r_data[7564];
                
                r_data[7566] <= r_data[7565];
                
                r_data[7567] <= r_data[7566];
                
                r_data[7568] <= r_data[7567];
                
                r_data[7569] <= r_data[7568];
                
                r_data[7570] <= r_data[7569];
                
                r_data[7571] <= r_data[7570];
                
                r_data[7572] <= r_data[7571];
                
                r_data[7573] <= r_data[7572];
                
                r_data[7574] <= r_data[7573];
                
                r_data[7575] <= r_data[7574];
                
                r_data[7576] <= r_data[7575];
                
                r_data[7577] <= r_data[7576];
                
                r_data[7578] <= r_data[7577];
                
                r_data[7579] <= r_data[7578];
                
                r_data[7580] <= r_data[7579];
                
                r_data[7581] <= r_data[7580];
                
                r_data[7582] <= r_data[7581];
                
                r_data[7583] <= r_data[7582];
                
                r_data[7584] <= r_data[7583];
                
                r_data[7585] <= r_data[7584];
                
                r_data[7586] <= r_data[7585];
                
                r_data[7587] <= r_data[7586];
                
                r_data[7588] <= r_data[7587];
                
                r_data[7589] <= r_data[7588];
                
                r_data[7590] <= r_data[7589];
                
                r_data[7591] <= r_data[7590];
                
                r_data[7592] <= r_data[7591];
                
                r_data[7593] <= r_data[7592];
                
                r_data[7594] <= r_data[7593];
                
                r_data[7595] <= r_data[7594];
                
                r_data[7596] <= r_data[7595];
                
                r_data[7597] <= r_data[7596];
                
                r_data[7598] <= r_data[7597];
                
                r_data[7599] <= r_data[7598];
                
                r_data[7600] <= r_data[7599];
                
                r_data[7601] <= r_data[7600];
                
                r_data[7602] <= r_data[7601];
                
                r_data[7603] <= r_data[7602];
                
                r_data[7604] <= r_data[7603];
                
                r_data[7605] <= r_data[7604];
                
                r_data[7606] <= r_data[7605];
                
                r_data[7607] <= r_data[7606];
                
                r_data[7608] <= r_data[7607];
                
                r_data[7609] <= r_data[7608];
                
                r_data[7610] <= r_data[7609];
                
                r_data[7611] <= r_data[7610];
                
                r_data[7612] <= r_data[7611];
                
                r_data[7613] <= r_data[7612];
                
                r_data[7614] <= r_data[7613];
                
                r_data[7615] <= r_data[7614];
                
                r_data[7616] <= r_data[7615];
                
                r_data[7617] <= r_data[7616];
                
                r_data[7618] <= r_data[7617];
                
                r_data[7619] <= r_data[7618];
                
                r_data[7620] <= r_data[7619];
                
                r_data[7621] <= r_data[7620];
                
                r_data[7622] <= r_data[7621];
                
                r_data[7623] <= r_data[7622];
                
                r_data[7624] <= r_data[7623];
                
                r_data[7625] <= r_data[7624];
                
                r_data[7626] <= r_data[7625];
                
                r_data[7627] <= r_data[7626];
                
                r_data[7628] <= r_data[7627];
                
                r_data[7629] <= r_data[7628];
                
                r_data[7630] <= r_data[7629];
                
                r_data[7631] <= r_data[7630];
                
                r_data[7632] <= r_data[7631];
                
                r_data[7633] <= r_data[7632];
                
                r_data[7634] <= r_data[7633];
                
                r_data[7635] <= r_data[7634];
                
                r_data[7636] <= r_data[7635];
                
                r_data[7637] <= r_data[7636];
                
                r_data[7638] <= r_data[7637];
                
                r_data[7639] <= r_data[7638];
                
                r_data[7640] <= r_data[7639];
                
                r_data[7641] <= r_data[7640];
                
                r_data[7642] <= r_data[7641];
                
                r_data[7643] <= r_data[7642];
                
                r_data[7644] <= r_data[7643];
                
                r_data[7645] <= r_data[7644];
                
                r_data[7646] <= r_data[7645];
                
                r_data[7647] <= r_data[7646];
                
                r_data[7648] <= r_data[7647];
                
                r_data[7649] <= r_data[7648];
                
                r_data[7650] <= r_data[7649];
                
                r_data[7651] <= r_data[7650];
                
                r_data[7652] <= r_data[7651];
                
                r_data[7653] <= r_data[7652];
                
                r_data[7654] <= r_data[7653];
                
                r_data[7655] <= r_data[7654];
                
                r_data[7656] <= r_data[7655];
                
                r_data[7657] <= r_data[7656];
                
                r_data[7658] <= r_data[7657];
                
                r_data[7659] <= r_data[7658];
                
                r_data[7660] <= r_data[7659];
                
                r_data[7661] <= r_data[7660];
                
                r_data[7662] <= r_data[7661];
                
                r_data[7663] <= r_data[7662];
                
                r_data[7664] <= r_data[7663];
                
                r_data[7665] <= r_data[7664];
                
                r_data[7666] <= r_data[7665];
                
                r_data[7667] <= r_data[7666];
                
                r_data[7668] <= r_data[7667];
                
                r_data[7669] <= r_data[7668];
                
                r_data[7670] <= r_data[7669];
                
                r_data[7671] <= r_data[7670];
                
                r_data[7672] <= r_data[7671];
                
                r_data[7673] <= r_data[7672];
                
                r_data[7674] <= r_data[7673];
                
                r_data[7675] <= r_data[7674];
                
                r_data[7676] <= r_data[7675];
                
                r_data[7677] <= r_data[7676];
                
                r_data[7678] <= r_data[7677];
                
                r_data[7679] <= r_data[7678];
                
                r_data[7680] <= r_data[7679];
                
                r_data[7681] <= r_data[7680];
                
                r_data[7682] <= r_data[7681];
                
                r_data[7683] <= r_data[7682];
                
                r_data[7684] <= r_data[7683];
                
                r_data[7685] <= r_data[7684];
                
                r_data[7686] <= r_data[7685];
                
                r_data[7687] <= r_data[7686];
                
                r_data[7688] <= r_data[7687];
                
                r_data[7689] <= r_data[7688];
                
                r_data[7690] <= r_data[7689];
                
                r_data[7691] <= r_data[7690];
                
                r_data[7692] <= r_data[7691];
                
                r_data[7693] <= r_data[7692];
                
                r_data[7694] <= r_data[7693];
                
                r_data[7695] <= r_data[7694];
                
                r_data[7696] <= r_data[7695];
                
                r_data[7697] <= r_data[7696];
                
                r_data[7698] <= r_data[7697];
                
                r_data[7699] <= r_data[7698];
                
                r_data[7700] <= r_data[7699];
                
                r_data[7701] <= r_data[7700];
                
                r_data[7702] <= r_data[7701];
                
                r_data[7703] <= r_data[7702];
                
                r_data[7704] <= r_data[7703];
                
                r_data[7705] <= r_data[7704];
                
                r_data[7706] <= r_data[7705];
                
                r_data[7707] <= r_data[7706];
                
                r_data[7708] <= r_data[7707];
                
                r_data[7709] <= r_data[7708];
                
                r_data[7710] <= r_data[7709];
                
                r_data[7711] <= r_data[7710];
                
                r_data[7712] <= r_data[7711];
                
                r_data[7713] <= r_data[7712];
                
                r_data[7714] <= r_data[7713];
                
                r_data[7715] <= r_data[7714];
                
                r_data[7716] <= r_data[7715];
                
                r_data[7717] <= r_data[7716];
                
                r_data[7718] <= r_data[7717];
                
                r_data[7719] <= r_data[7718];
                
                r_data[7720] <= r_data[7719];
                
                r_data[7721] <= r_data[7720];
                
                r_data[7722] <= r_data[7721];
                
                r_data[7723] <= r_data[7722];
                
                r_data[7724] <= r_data[7723];
                
                r_data[7725] <= r_data[7724];
                
                r_data[7726] <= r_data[7725];
                
                r_data[7727] <= r_data[7726];
                
                r_data[7728] <= r_data[7727];
                
                r_data[7729] <= r_data[7728];
                
                r_data[7730] <= r_data[7729];
                
                r_data[7731] <= r_data[7730];
                
                r_data[7732] <= r_data[7731];
                
                r_data[7733] <= r_data[7732];
                
                r_data[7734] <= r_data[7733];
                
                r_data[7735] <= r_data[7734];
                
                r_data[7736] <= r_data[7735];
                
                r_data[7737] <= r_data[7736];
                
                r_data[7738] <= r_data[7737];
                
                r_data[7739] <= r_data[7738];
                
                r_data[7740] <= r_data[7739];
                
                r_data[7741] <= r_data[7740];
                
                r_data[7742] <= r_data[7741];
                
                r_data[7743] <= r_data[7742];
                
                r_data[7744] <= r_data[7743];
                
                r_data[7745] <= r_data[7744];
                
                r_data[7746] <= r_data[7745];
                
                r_data[7747] <= r_data[7746];
                
                r_data[7748] <= r_data[7747];
                
                r_data[7749] <= r_data[7748];
                
                r_data[7750] <= r_data[7749];
                
                r_data[7751] <= r_data[7750];
                
                r_data[7752] <= r_data[7751];
                
                r_data[7753] <= r_data[7752];
                
                r_data[7754] <= r_data[7753];
                
                r_data[7755] <= r_data[7754];
                
                r_data[7756] <= r_data[7755];
                
                r_data[7757] <= r_data[7756];
                
                r_data[7758] <= r_data[7757];
                
                r_data[7759] <= r_data[7758];
                
                r_data[7760] <= r_data[7759];
                
                r_data[7761] <= r_data[7760];
                
                r_data[7762] <= r_data[7761];
                
                r_data[7763] <= r_data[7762];
                
                r_data[7764] <= r_data[7763];
                
                r_data[7765] <= r_data[7764];
                
                r_data[7766] <= r_data[7765];
                
                r_data[7767] <= r_data[7766];
                
                r_data[7768] <= r_data[7767];
                
                r_data[7769] <= r_data[7768];
                
                r_data[7770] <= r_data[7769];
                
                r_data[7771] <= r_data[7770];
                
                r_data[7772] <= r_data[7771];
                
                r_data[7773] <= r_data[7772];
                
                r_data[7774] <= r_data[7773];
                
                r_data[7775] <= r_data[7774];
                
                r_data[7776] <= r_data[7775];
                
                r_data[7777] <= r_data[7776];
                
                r_data[7778] <= r_data[7777];
                
                r_data[7779] <= r_data[7778];
                
                r_data[7780] <= r_data[7779];
                
                r_data[7781] <= r_data[7780];
                
                r_data[7782] <= r_data[7781];
                
                r_data[7783] <= r_data[7782];
                
                r_data[7784] <= r_data[7783];
                
                r_data[7785] <= r_data[7784];
                
                r_data[7786] <= r_data[7785];
                
                r_data[7787] <= r_data[7786];
                
                r_data[7788] <= r_data[7787];
                
                r_data[7789] <= r_data[7788];
                
                r_data[7790] <= r_data[7789];
                
                r_data[7791] <= r_data[7790];
                
                r_data[7792] <= r_data[7791];
                
                r_data[7793] <= r_data[7792];
                
                r_data[7794] <= r_data[7793];
                
                r_data[7795] <= r_data[7794];
                
                r_data[7796] <= r_data[7795];
                
                r_data[7797] <= r_data[7796];
                
                r_data[7798] <= r_data[7797];
                
                r_data[7799] <= r_data[7798];
                
                r_data[7800] <= r_data[7799];
                
                r_data[7801] <= r_data[7800];
                
                r_data[7802] <= r_data[7801];
                
                r_data[7803] <= r_data[7802];
                
                r_data[7804] <= r_data[7803];
                
                r_data[7805] <= r_data[7804];
                
                r_data[7806] <= r_data[7805];
                
                r_data[7807] <= r_data[7806];
                
                r_data[7808] <= r_data[7807];
                
                r_data[7809] <= r_data[7808];
                
                r_data[7810] <= r_data[7809];
                
                r_data[7811] <= r_data[7810];
                
                r_data[7812] <= r_data[7811];
                
                r_data[7813] <= r_data[7812];
                
                r_data[7814] <= r_data[7813];
                
                r_data[7815] <= r_data[7814];
                
                r_data[7816] <= r_data[7815];
                
                r_data[7817] <= r_data[7816];
                
                r_data[7818] <= r_data[7817];
                
                r_data[7819] <= r_data[7818];
                
                r_data[7820] <= r_data[7819];
                
                r_data[7821] <= r_data[7820];
                
                r_data[7822] <= r_data[7821];
                
                r_data[7823] <= r_data[7822];
                
                r_data[7824] <= r_data[7823];
                
                r_data[7825] <= r_data[7824];
                
                r_data[7826] <= r_data[7825];
                
                r_data[7827] <= r_data[7826];
                
                r_data[7828] <= r_data[7827];
                
                r_data[7829] <= r_data[7828];
                
                r_data[7830] <= r_data[7829];
                
                r_data[7831] <= r_data[7830];
                
                r_data[7832] <= r_data[7831];
                
                r_data[7833] <= r_data[7832];
                
                r_data[7834] <= r_data[7833];
                
                r_data[7835] <= r_data[7834];
                
                r_data[7836] <= r_data[7835];
                
                r_data[7837] <= r_data[7836];
                
                r_data[7838] <= r_data[7837];
                
                r_data[7839] <= r_data[7838];
                
                r_data[7840] <= r_data[7839];
                
                r_data[7841] <= r_data[7840];
                
                r_data[7842] <= r_data[7841];
                
                r_data[7843] <= r_data[7842];
                
                r_data[7844] <= r_data[7843];
                
                r_data[7845] <= r_data[7844];
                
                r_data[7846] <= r_data[7845];
                
                r_data[7847] <= r_data[7846];
                
                r_data[7848] <= r_data[7847];
                
                r_data[7849] <= r_data[7848];
                
                r_data[7850] <= r_data[7849];
                
                r_data[7851] <= r_data[7850];
                
                r_data[7852] <= r_data[7851];
                
                r_data[7853] <= r_data[7852];
                
                r_data[7854] <= r_data[7853];
                
                r_data[7855] <= r_data[7854];
                
                r_data[7856] <= r_data[7855];
                
                r_data[7857] <= r_data[7856];
                
                r_data[7858] <= r_data[7857];
                
                r_data[7859] <= r_data[7858];
                
                r_data[7860] <= r_data[7859];
                
                r_data[7861] <= r_data[7860];
                
                r_data[7862] <= r_data[7861];
                
                r_data[7863] <= r_data[7862];
                
                r_data[7864] <= r_data[7863];
                
                r_data[7865] <= r_data[7864];
                
                r_data[7866] <= r_data[7865];
                
                r_data[7867] <= r_data[7866];
                
                r_data[7868] <= r_data[7867];
                
                r_data[7869] <= r_data[7868];
                
                r_data[7870] <= r_data[7869];
                
                r_data[7871] <= r_data[7870];
                
                r_data[7872] <= r_data[7871];
                
                r_data[7873] <= r_data[7872];
                
                r_data[7874] <= r_data[7873];
                
                r_data[7875] <= r_data[7874];
                
                r_data[7876] <= r_data[7875];
                
                r_data[7877] <= r_data[7876];
                
                r_data[7878] <= r_data[7877];
                
                r_data[7879] <= r_data[7878];
                
                r_data[7880] <= r_data[7879];
                
                r_data[7881] <= r_data[7880];
                
                r_data[7882] <= r_data[7881];
                
                r_data[7883] <= r_data[7882];
                
                r_data[7884] <= r_data[7883];
                
                r_data[7885] <= r_data[7884];
                
                r_data[7886] <= r_data[7885];
                
                r_data[7887] <= r_data[7886];
                
                r_data[7888] <= r_data[7887];
                
                r_data[7889] <= r_data[7888];
                
                r_data[7890] <= r_data[7889];
                
                r_data[7891] <= r_data[7890];
                
                r_data[7892] <= r_data[7891];
                
                r_data[7893] <= r_data[7892];
                
                r_data[7894] <= r_data[7893];
                
                r_data[7895] <= r_data[7894];
                
                r_data[7896] <= r_data[7895];
                
                r_data[7897] <= r_data[7896];
                
                r_data[7898] <= r_data[7897];
                
                r_data[7899] <= r_data[7898];
                
                r_data[7900] <= r_data[7899];
                
                r_data[7901] <= r_data[7900];
                
                r_data[7902] <= r_data[7901];
                
                r_data[7903] <= r_data[7902];
                
                r_data[7904] <= r_data[7903];
                
                r_data[7905] <= r_data[7904];
                
                r_data[7906] <= r_data[7905];
                
                r_data[7907] <= r_data[7906];
                
                r_data[7908] <= r_data[7907];
                
                r_data[7909] <= r_data[7908];
                
                r_data[7910] <= r_data[7909];
                
                r_data[7911] <= r_data[7910];
                
                r_data[7912] <= r_data[7911];
                
                r_data[7913] <= r_data[7912];
                
                r_data[7914] <= r_data[7913];
                
                r_data[7915] <= r_data[7914];
                
                r_data[7916] <= r_data[7915];
                
                r_data[7917] <= r_data[7916];
                
                r_data[7918] <= r_data[7917];
                
                r_data[7919] <= r_data[7918];
                
                r_data[7920] <= r_data[7919];
                
                r_data[7921] <= r_data[7920];
                
                r_data[7922] <= r_data[7921];
                
                r_data[7923] <= r_data[7922];
                
                r_data[7924] <= r_data[7923];
                
                r_data[7925] <= r_data[7924];
                
                r_data[7926] <= r_data[7925];
                
                r_data[7927] <= r_data[7926];
                
                r_data[7928] <= r_data[7927];
                
                r_data[7929] <= r_data[7928];
                
                r_data[7930] <= r_data[7929];
                
                r_data[7931] <= r_data[7930];
                
                r_data[7932] <= r_data[7931];
                
                r_data[7933] <= r_data[7932];
                
                r_data[7934] <= r_data[7933];
                
                r_data[7935] <= r_data[7934];
                
                r_data[7936] <= r_data[7935];
                
                r_data[7937] <= r_data[7936];
                
                r_data[7938] <= r_data[7937];
                
                r_data[7939] <= r_data[7938];
                
                r_data[7940] <= r_data[7939];
                
                r_data[7941] <= r_data[7940];
                
                r_data[7942] <= r_data[7941];
                
                r_data[7943] <= r_data[7942];
                
                r_data[7944] <= r_data[7943];
                
                r_data[7945] <= r_data[7944];
                
                r_data[7946] <= r_data[7945];
                
                r_data[7947] <= r_data[7946];
                
                r_data[7948] <= r_data[7947];
                
                r_data[7949] <= r_data[7948];
                
                r_data[7950] <= r_data[7949];
                
                r_data[7951] <= r_data[7950];
                
                r_data[7952] <= r_data[7951];
                
                r_data[7953] <= r_data[7952];
                
                r_data[7954] <= r_data[7953];
                
                r_data[7955] <= r_data[7954];
                
                r_data[7956] <= r_data[7955];
                
                r_data[7957] <= r_data[7956];
                
                r_data[7958] <= r_data[7957];
                
                r_data[7959] <= r_data[7958];
                
                r_data[7960] <= r_data[7959];
                
                r_data[7961] <= r_data[7960];
                
                r_data[7962] <= r_data[7961];
                
                r_data[7963] <= r_data[7962];
                
                r_data[7964] <= r_data[7963];
                
                r_data[7965] <= r_data[7964];
                
                r_data[7966] <= r_data[7965];
                
                r_data[7967] <= r_data[7966];
                
                r_data[7968] <= r_data[7967];
                
                r_data[7969] <= r_data[7968];
                
                r_data[7970] <= r_data[7969];
                
                r_data[7971] <= r_data[7970];
                
                r_data[7972] <= r_data[7971];
                
                r_data[7973] <= r_data[7972];
                
                r_data[7974] <= r_data[7973];
                
                r_data[7975] <= r_data[7974];
                
                r_data[7976] <= r_data[7975];
                
                r_data[7977] <= r_data[7976];
                
                r_data[7978] <= r_data[7977];
                
                r_data[7979] <= r_data[7978];
                
                r_data[7980] <= r_data[7979];
                
                r_data[7981] <= r_data[7980];
                
                r_data[7982] <= r_data[7981];
                
                r_data[7983] <= r_data[7982];
                
                r_data[7984] <= r_data[7983];
                
                r_data[7985] <= r_data[7984];
                
                r_data[7986] <= r_data[7985];
                
                r_data[7987] <= r_data[7986];
                
                r_data[7988] <= r_data[7987];
                
                r_data[7989] <= r_data[7988];
                
                r_data[7990] <= r_data[7989];
                
                r_data[7991] <= r_data[7990];
                
                r_data[7992] <= r_data[7991];
                
                r_data[7993] <= r_data[7992];
                
                r_data[7994] <= r_data[7993];
                
                r_data[7995] <= r_data[7994];
                
                r_data[7996] <= r_data[7995];
                
                r_data[7997] <= r_data[7996];
                
                r_data[7998] <= r_data[7997];
                
                r_data[7999] <= r_data[7998];
                
                r_data[8000] <= r_data[7999];
                
                r_data[8001] <= r_data[8000];
                
                r_data[8002] <= r_data[8001];
                
                r_data[8003] <= r_data[8002];
                
                r_data[8004] <= r_data[8003];
                
                r_data[8005] <= r_data[8004];
                
                r_data[8006] <= r_data[8005];
                
                r_data[8007] <= r_data[8006];
                
                r_data[8008] <= r_data[8007];
                
                r_data[8009] <= r_data[8008];
                
                r_data[8010] <= r_data[8009];
                
                r_data[8011] <= r_data[8010];
                
                r_data[8012] <= r_data[8011];
                
                r_data[8013] <= r_data[8012];
                
                r_data[8014] <= r_data[8013];
                
                r_data[8015] <= r_data[8014];
                
                r_data[8016] <= r_data[8015];
                
                r_data[8017] <= r_data[8016];
                
                r_data[8018] <= r_data[8017];
                
                r_data[8019] <= r_data[8018];
                
                r_data[8020] <= r_data[8019];
                
                r_data[8021] <= r_data[8020];
                
                r_data[8022] <= r_data[8021];
                
                r_data[8023] <= r_data[8022];
                
                r_data[8024] <= r_data[8023];
                
                r_data[8025] <= r_data[8024];
                
                r_data[8026] <= r_data[8025];
                
                r_data[8027] <= r_data[8026];
                
                r_data[8028] <= r_data[8027];
                
                r_data[8029] <= r_data[8028];
                
                r_data[8030] <= r_data[8029];
                
                r_data[8031] <= r_data[8030];
                
                r_data[8032] <= r_data[8031];
                
                r_data[8033] <= r_data[8032];
                
                r_data[8034] <= r_data[8033];
                
                r_data[8035] <= r_data[8034];
                
                r_data[8036] <= r_data[8035];
                
                r_data[8037] <= r_data[8036];
                
                r_data[8038] <= r_data[8037];
                
                r_data[8039] <= r_data[8038];
                
                r_data[8040] <= r_data[8039];
                
                r_data[8041] <= r_data[8040];
                
                r_data[8042] <= r_data[8041];
                
                r_data[8043] <= r_data[8042];
                
                r_data[8044] <= r_data[8043];
                
                r_data[8045] <= r_data[8044];
                
                r_data[8046] <= r_data[8045];
                
                r_data[8047] <= r_data[8046];
                
                r_data[8048] <= r_data[8047];
                
                r_data[8049] <= r_data[8048];
                
                r_data[8050] <= r_data[8049];
                
                r_data[8051] <= r_data[8050];
                
                r_data[8052] <= r_data[8051];
                
                r_data[8053] <= r_data[8052];
                
                r_data[8054] <= r_data[8053];
                
                r_data[8055] <= r_data[8054];
                
                r_data[8056] <= r_data[8055];
                
                r_data[8057] <= r_data[8056];
                
                r_data[8058] <= r_data[8057];
                
                r_data[8059] <= r_data[8058];
                
                r_data[8060] <= r_data[8059];
                
                r_data[8061] <= r_data[8060];
                
                r_data[8062] <= r_data[8061];
                
                r_data[8063] <= r_data[8062];
                
                r_data[8064] <= r_data[8063];
                
                r_data[8065] <= r_data[8064];
                
                r_data[8066] <= r_data[8065];
                
                r_data[8067] <= r_data[8066];
                
                r_data[8068] <= r_data[8067];
                
                r_data[8069] <= r_data[8068];
                
                r_data[8070] <= r_data[8069];
                
                r_data[8071] <= r_data[8070];
                
                r_data[8072] <= r_data[8071];
                
                r_data[8073] <= r_data[8072];
                
                r_data[8074] <= r_data[8073];
                
                r_data[8075] <= r_data[8074];
                
                r_data[8076] <= r_data[8075];
                
                r_data[8077] <= r_data[8076];
                
                r_data[8078] <= r_data[8077];
                
                r_data[8079] <= r_data[8078];
                
                r_data[8080] <= r_data[8079];
                
                r_data[8081] <= r_data[8080];
                
                r_data[8082] <= r_data[8081];
                
                r_data[8083] <= r_data[8082];
                
                r_data[8084] <= r_data[8083];
                
                r_data[8085] <= r_data[8084];
                
                r_data[8086] <= r_data[8085];
                
                r_data[8087] <= r_data[8086];
                
                r_data[8088] <= r_data[8087];
                
                r_data[8089] <= r_data[8088];
                
                r_data[8090] <= r_data[8089];
                
                r_data[8091] <= r_data[8090];
                
                r_data[8092] <= r_data[8091];
                
                r_data[8093] <= r_data[8092];
                
                r_data[8094] <= r_data[8093];
                
                r_data[8095] <= r_data[8094];
                
                r_data[8096] <= r_data[8095];
                
                r_data[8097] <= r_data[8096];
                
                r_data[8098] <= r_data[8097];
                
                r_data[8099] <= r_data[8098];
                
                r_data[8100] <= r_data[8099];
                
                r_data[8101] <= r_data[8100];
                
                r_data[8102] <= r_data[8101];
                
                r_data[8103] <= r_data[8102];
                
                r_data[8104] <= r_data[8103];
                
                r_data[8105] <= r_data[8104];
                
                r_data[8106] <= r_data[8105];
                
                r_data[8107] <= r_data[8106];
                
                r_data[8108] <= r_data[8107];
                
                r_data[8109] <= r_data[8108];
                
                r_data[8110] <= r_data[8109];
                
                r_data[8111] <= r_data[8110];
                
                r_data[8112] <= r_data[8111];
                
                r_data[8113] <= r_data[8112];
                
                r_data[8114] <= r_data[8113];
                
                r_data[8115] <= r_data[8114];
                
                r_data[8116] <= r_data[8115];
                
                r_data[8117] <= r_data[8116];
                
                r_data[8118] <= r_data[8117];
                
                r_data[8119] <= r_data[8118];
                
                r_data[8120] <= r_data[8119];
                
                r_data[8121] <= r_data[8120];
                
                r_data[8122] <= r_data[8121];
                
                r_data[8123] <= r_data[8122];
                
                r_data[8124] <= r_data[8123];
                
                r_data[8125] <= r_data[8124];
                
                r_data[8126] <= r_data[8125];
                
                r_data[8127] <= r_data[8126];
                
                r_data[8128] <= r_data[8127];
                
                r_data[8129] <= r_data[8128];
                
                r_data[8130] <= r_data[8129];
                
                r_data[8131] <= r_data[8130];
                
                r_data[8132] <= r_data[8131];
                
                r_data[8133] <= r_data[8132];
                
                r_data[8134] <= r_data[8133];
                
                r_data[8135] <= r_data[8134];
                
                r_data[8136] <= r_data[8135];
                
                r_data[8137] <= r_data[8136];
                
                r_data[8138] <= r_data[8137];
                
                r_data[8139] <= r_data[8138];
                
                r_data[8140] <= r_data[8139];
                
                r_data[8141] <= r_data[8140];
                
                r_data[8142] <= r_data[8141];
                
                r_data[8143] <= r_data[8142];
                
                r_data[8144] <= r_data[8143];
                
                r_data[8145] <= r_data[8144];
                
                r_data[8146] <= r_data[8145];
                
                r_data[8147] <= r_data[8146];
                
                r_data[8148] <= r_data[8147];
                
                r_data[8149] <= r_data[8148];
                
                r_data[8150] <= r_data[8149];
                
                r_data[8151] <= r_data[8150];
                
                r_data[8152] <= r_data[8151];
                
                r_data[8153] <= r_data[8152];
                
                r_data[8154] <= r_data[8153];
                
                r_data[8155] <= r_data[8154];
                
                r_data[8156] <= r_data[8155];
                
                r_data[8157] <= r_data[8156];
                
                r_data[8158] <= r_data[8157];
                
                r_data[8159] <= r_data[8158];
                
                r_data[8160] <= r_data[8159];
                
                r_data[8161] <= r_data[8160];
                
                r_data[8162] <= r_data[8161];
                
                r_data[8163] <= r_data[8162];
                
                r_data[8164] <= r_data[8163];
                
                r_data[8165] <= r_data[8164];
                
                r_data[8166] <= r_data[8165];
                
                r_data[8167] <= r_data[8166];
                
                r_data[8168] <= r_data[8167];
                
                r_data[8169] <= r_data[8168];
                
                r_data[8170] <= r_data[8169];
                
                r_data[8171] <= r_data[8170];
                
                r_data[8172] <= r_data[8171];
                
                r_data[8173] <= r_data[8172];
                
                r_data[8174] <= r_data[8173];
                
                r_data[8175] <= r_data[8174];
                
                r_data[8176] <= r_data[8175];
                
                r_data[8177] <= r_data[8176];
                
                r_data[8178] <= r_data[8177];
                
                r_data[8179] <= r_data[8178];
                
                r_data[8180] <= r_data[8179];
                
                r_data[8181] <= r_data[8180];
                
                r_data[8182] <= r_data[8181];
                
                r_data[8183] <= r_data[8182];
                
                r_data[8184] <= r_data[8183];
                
                r_data[8185] <= r_data[8184];
                
                r_data[8186] <= r_data[8185];
                
                r_data[8187] <= r_data[8186];
                
                r_data[8188] <= r_data[8187];
                
                r_data[8189] <= r_data[8188];
                
                r_data[8190] <= r_data[8189];
                
                r_data[8191] <= r_data[8190];
                
                r_data[8192] <= r_data[8191];
                
                r_data[8193] <= r_data[8192];
                
                r_data[8194] <= r_data[8193];
                
                r_data[8195] <= r_data[8194];
                
                r_data[8196] <= r_data[8195];
                
                r_data[8197] <= r_data[8196];
                
                r_data[8198] <= r_data[8197];
                
                r_data[8199] <= r_data[8198];
                
                r_data[8200] <= r_data[8199];
                
                r_data[8201] <= r_data[8200];
                
                r_data[8202] <= r_data[8201];
                
                r_data[8203] <= r_data[8202];
                
                r_data[8204] <= r_data[8203];
                
                r_data[8205] <= r_data[8204];
                
                r_data[8206] <= r_data[8205];
                
                r_data[8207] <= r_data[8206];
                
                r_data[8208] <= r_data[8207];
                
                r_data[8209] <= r_data[8208];
                
                r_data[8210] <= r_data[8209];
                
                r_data[8211] <= r_data[8210];
                
                r_data[8212] <= r_data[8211];
                
                r_data[8213] <= r_data[8212];
                
                r_data[8214] <= r_data[8213];
                
                r_data[8215] <= r_data[8214];
                
                r_data[8216] <= r_data[8215];
                
                r_data[8217] <= r_data[8216];
                
                r_data[8218] <= r_data[8217];
                
                r_data[8219] <= r_data[8218];
                
                r_data[8220] <= r_data[8219];
                
                r_data[8221] <= r_data[8220];
                
                r_data[8222] <= r_data[8221];
                
                r_data[8223] <= r_data[8222];
                
                r_data[8224] <= r_data[8223];
                
                r_data[8225] <= r_data[8224];
                
                r_data[8226] <= r_data[8225];
                
                r_data[8227] <= r_data[8226];
                
                r_data[8228] <= r_data[8227];
                
                r_data[8229] <= r_data[8228];
                
                r_data[8230] <= r_data[8229];
                
                r_data[8231] <= r_data[8230];
                
                r_data[8232] <= r_data[8231];
                
                r_data[8233] <= r_data[8232];
                
                r_data[8234] <= r_data[8233];
                
                r_data[8235] <= r_data[8234];
                
                r_data[8236] <= r_data[8235];
                
                r_data[8237] <= r_data[8236];
                
                r_data[8238] <= r_data[8237];
                
                r_data[8239] <= r_data[8238];
                
                r_data[8240] <= r_data[8239];
                
                r_data[8241] <= r_data[8240];
                
                r_data[8242] <= r_data[8241];
                
                r_data[8243] <= r_data[8242];
                
                r_data[8244] <= r_data[8243];
                
                r_data[8245] <= r_data[8244];
                
                r_data[8246] <= r_data[8245];
                
                r_data[8247] <= r_data[8246];
                
                r_data[8248] <= r_data[8247];
                
                r_data[8249] <= r_data[8248];
                
                r_data[8250] <= r_data[8249];
                
                r_data[8251] <= r_data[8250];
                
                r_data[8252] <= r_data[8251];
                
                r_data[8253] <= r_data[8252];
                
                r_data[8254] <= r_data[8253];
                
                r_data[8255] <= r_data[8254];
                
                r_data[8256] <= r_data[8255];
                
                r_data[8257] <= r_data[8256];
                
                r_data[8258] <= r_data[8257];
                
                r_data[8259] <= r_data[8258];
                
                r_data[8260] <= r_data[8259];
                
                r_data[8261] <= r_data[8260];
                
                r_data[8262] <= r_data[8261];
                
                r_data[8263] <= r_data[8262];
                
                r_data[8264] <= r_data[8263];
                
                r_data[8265] <= r_data[8264];
                
                r_data[8266] <= r_data[8265];
                
                r_data[8267] <= r_data[8266];
                
                r_data[8268] <= r_data[8267];
                
                r_data[8269] <= r_data[8268];
                
                r_data[8270] <= r_data[8269];
                
                r_data[8271] <= r_data[8270];
                
                r_data[8272] <= r_data[8271];
                
                r_data[8273] <= r_data[8272];
                
                r_data[8274] <= r_data[8273];
                
                r_data[8275] <= r_data[8274];
                
                r_data[8276] <= r_data[8275];
                
                r_data[8277] <= r_data[8276];
                
                r_data[8278] <= r_data[8277];
                
                r_data[8279] <= r_data[8278];
                
                r_data[8280] <= r_data[8279];
                
                r_data[8281] <= r_data[8280];
                
                r_data[8282] <= r_data[8281];
                
                r_data[8283] <= r_data[8282];
                
                r_data[8284] <= r_data[8283];
                
                r_data[8285] <= r_data[8284];
                
                r_data[8286] <= r_data[8285];
                
                r_data[8287] <= r_data[8286];
                
                r_data[8288] <= r_data[8287];
                
                r_data[8289] <= r_data[8288];
                
                r_data[8290] <= r_data[8289];
                
                r_data[8291] <= r_data[8290];
                
                r_data[8292] <= r_data[8291];
                
                r_data[8293] <= r_data[8292];
                
                r_data[8294] <= r_data[8293];
                
                r_data[8295] <= r_data[8294];
                
                r_data[8296] <= r_data[8295];
                
                r_data[8297] <= r_data[8296];
                
                r_data[8298] <= r_data[8297];
                
                r_data[8299] <= r_data[8298];
                
                r_data[8300] <= r_data[8299];
                
                r_data[8301] <= r_data[8300];
                
                r_data[8302] <= r_data[8301];
                
                r_data[8303] <= r_data[8302];
                
                r_data[8304] <= r_data[8303];
                
                r_data[8305] <= r_data[8304];
                
                r_data[8306] <= r_data[8305];
                
                r_data[8307] <= r_data[8306];
                
                r_data[8308] <= r_data[8307];
                
                r_data[8309] <= r_data[8308];
                
                r_data[8310] <= r_data[8309];
                
                r_data[8311] <= r_data[8310];
                
                r_data[8312] <= r_data[8311];
                
                r_data[8313] <= r_data[8312];
                
                r_data[8314] <= r_data[8313];
                
                r_data[8315] <= r_data[8314];
                
                r_data[8316] <= r_data[8315];
                
                r_data[8317] <= r_data[8316];
                
                r_data[8318] <= r_data[8317];
                
                r_data[8319] <= r_data[8318];
                
                r_data[8320] <= r_data[8319];
                
                r_data[8321] <= r_data[8320];
                
                r_data[8322] <= r_data[8321];
                
                r_data[8323] <= r_data[8322];
                
                r_data[8324] <= r_data[8323];
                
                r_data[8325] <= r_data[8324];
                
                r_data[8326] <= r_data[8325];
                
                r_data[8327] <= r_data[8326];
                
                r_data[8328] <= r_data[8327];
                
                r_data[8329] <= r_data[8328];
                
                r_data[8330] <= r_data[8329];
                
                r_data[8331] <= r_data[8330];
                
                r_data[8332] <= r_data[8331];
                
                r_data[8333] <= r_data[8332];
                
                r_data[8334] <= r_data[8333];
                
                r_data[8335] <= r_data[8334];
                
                r_data[8336] <= r_data[8335];
                
                r_data[8337] <= r_data[8336];
                
                r_data[8338] <= r_data[8337];
                
                r_data[8339] <= r_data[8338];
                
                r_data[8340] <= r_data[8339];
                
                r_data[8341] <= r_data[8340];
                
                r_data[8342] <= r_data[8341];
                
                r_data[8343] <= r_data[8342];
                
                r_data[8344] <= r_data[8343];
                
                r_data[8345] <= r_data[8344];
                
                r_data[8346] <= r_data[8345];
                
                r_data[8347] <= r_data[8346];
                
                r_data[8348] <= r_data[8347];
                
                r_data[8349] <= r_data[8348];
                
                r_data[8350] <= r_data[8349];
                
                r_data[8351] <= r_data[8350];
                
                r_data[8352] <= r_data[8351];
                
                r_data[8353] <= r_data[8352];
                
                r_data[8354] <= r_data[8353];
                
                r_data[8355] <= r_data[8354];
                
                r_data[8356] <= r_data[8355];
                
                r_data[8357] <= r_data[8356];
                
                r_data[8358] <= r_data[8357];
                
                r_data[8359] <= r_data[8358];
                
                r_data[8360] <= r_data[8359];
                
                r_data[8361] <= r_data[8360];
                
                r_data[8362] <= r_data[8361];
                
                r_data[8363] <= r_data[8362];
                
                r_data[8364] <= r_data[8363];
                
                r_data[8365] <= r_data[8364];
                
                r_data[8366] <= r_data[8365];
                
                r_data[8367] <= r_data[8366];
                
                r_data[8368] <= r_data[8367];
                
                r_data[8369] <= r_data[8368];
                
                r_data[8370] <= r_data[8369];
                
                r_data[8371] <= r_data[8370];
                
                r_data[8372] <= r_data[8371];
                
                r_data[8373] <= r_data[8372];
                
                r_data[8374] <= r_data[8373];
                
                r_data[8375] <= r_data[8374];
                
                r_data[8376] <= r_data[8375];
                
                r_data[8377] <= r_data[8376];
                
                r_data[8378] <= r_data[8377];
                
                r_data[8379] <= r_data[8378];
                
                r_data[8380] <= r_data[8379];
                
                r_data[8381] <= r_data[8380];
                
                r_data[8382] <= r_data[8381];
                
                r_data[8383] <= r_data[8382];
                
                r_data[8384] <= r_data[8383];
                
                r_data[8385] <= r_data[8384];
                
                r_data[8386] <= r_data[8385];
                
                r_data[8387] <= r_data[8386];
                
                r_data[8388] <= r_data[8387];
                
                r_data[8389] <= r_data[8388];
                
                r_data[8390] <= r_data[8389];
                
                r_data[8391] <= r_data[8390];
                
                r_data[8392] <= r_data[8391];
                
                r_data[8393] <= r_data[8392];
                
                r_data[8394] <= r_data[8393];
                
                r_data[8395] <= r_data[8394];
                
                r_data[8396] <= r_data[8395];
                
                r_data[8397] <= r_data[8396];
                
                r_data[8398] <= r_data[8397];
                
                r_data[8399] <= r_data[8398];
                
                r_data[8400] <= r_data[8399];
                
                r_data[8401] <= r_data[8400];
                
                r_data[8402] <= r_data[8401];
                
                r_data[8403] <= r_data[8402];
                
                r_data[8404] <= r_data[8403];
                
                r_data[8405] <= r_data[8404];
                
                r_data[8406] <= r_data[8405];
                
                r_data[8407] <= r_data[8406];
                
                r_data[8408] <= r_data[8407];
                
                r_data[8409] <= r_data[8408];
                
                r_data[8410] <= r_data[8409];
                
                r_data[8411] <= r_data[8410];
                
                r_data[8412] <= r_data[8411];
                
                r_data[8413] <= r_data[8412];
                
                r_data[8414] <= r_data[8413];
                
                r_data[8415] <= r_data[8414];
                
                r_data[8416] <= r_data[8415];
                
                r_data[8417] <= r_data[8416];
                
                r_data[8418] <= r_data[8417];
                
                r_data[8419] <= r_data[8418];
                
                r_data[8420] <= r_data[8419];
                
                r_data[8421] <= r_data[8420];
                
                r_data[8422] <= r_data[8421];
                
                r_data[8423] <= r_data[8422];
                
                r_data[8424] <= r_data[8423];
                
                r_data[8425] <= r_data[8424];
                
                r_data[8426] <= r_data[8425];
                
                r_data[8427] <= r_data[8426];
                
                r_data[8428] <= r_data[8427];
                
                r_data[8429] <= r_data[8428];
                
                r_data[8430] <= r_data[8429];
                
                r_data[8431] <= r_data[8430];
                
                r_data[8432] <= r_data[8431];
                
                r_data[8433] <= r_data[8432];
                
                r_data[8434] <= r_data[8433];
                
                r_data[8435] <= r_data[8434];
                
                r_data[8436] <= r_data[8435];
                
                r_data[8437] <= r_data[8436];
                
                r_data[8438] <= r_data[8437];
                
                r_data[8439] <= r_data[8438];
                
                r_data[8440] <= r_data[8439];
                
                r_data[8441] <= r_data[8440];
                
                r_data[8442] <= r_data[8441];
                
                r_data[8443] <= r_data[8442];
                
                r_data[8444] <= r_data[8443];
                
                r_data[8445] <= r_data[8444];
                
                r_data[8446] <= r_data[8445];
                
                r_data[8447] <= r_data[8446];
                
                r_data[8448] <= r_data[8447];
                
                r_data[8449] <= r_data[8448];
                
                r_data[8450] <= r_data[8449];
                
                r_data[8451] <= r_data[8450];
                
                r_data[8452] <= r_data[8451];
                
                r_data[8453] <= r_data[8452];
                
                r_data[8454] <= r_data[8453];
                
                r_data[8455] <= r_data[8454];
                
                r_data[8456] <= r_data[8455];
                
                r_data[8457] <= r_data[8456];
                
                r_data[8458] <= r_data[8457];
                
                r_data[8459] <= r_data[8458];
                
                r_data[8460] <= r_data[8459];
                
                r_data[8461] <= r_data[8460];
                
                r_data[8462] <= r_data[8461];
                
                r_data[8463] <= r_data[8462];
                
                r_data[8464] <= r_data[8463];
                
                r_data[8465] <= r_data[8464];
                
                r_data[8466] <= r_data[8465];
                
                r_data[8467] <= r_data[8466];
                
                r_data[8468] <= r_data[8467];
                
                r_data[8469] <= r_data[8468];
                
                r_data[8470] <= r_data[8469];
                
                r_data[8471] <= r_data[8470];
                
                r_data[8472] <= r_data[8471];
                
                r_data[8473] <= r_data[8472];
                
                r_data[8474] <= r_data[8473];
                
                r_data[8475] <= r_data[8474];
                
                r_data[8476] <= r_data[8475];
                
                r_data[8477] <= r_data[8476];
                
                r_data[8478] <= r_data[8477];
                
                r_data[8479] <= r_data[8478];
                
                r_data[8480] <= r_data[8479];
                
                r_data[8481] <= r_data[8480];
                
                r_data[8482] <= r_data[8481];
                
                r_data[8483] <= r_data[8482];
                
                r_data[8484] <= r_data[8483];
                
                r_data[8485] <= r_data[8484];
                
                r_data[8486] <= r_data[8485];
                
                r_data[8487] <= r_data[8486];
                
                r_data[8488] <= r_data[8487];
                
                r_data[8489] <= r_data[8488];
                
                r_data[8490] <= r_data[8489];
                
                r_data[8491] <= r_data[8490];
                
                r_data[8492] <= r_data[8491];
                
                r_data[8493] <= r_data[8492];
                
                r_data[8494] <= r_data[8493];
                
                r_data[8495] <= r_data[8494];
                
                r_data[8496] <= r_data[8495];
                
                r_data[8497] <= r_data[8496];
                
                r_data[8498] <= r_data[8497];
                
                r_data[8499] <= r_data[8498];
                
                r_data[8500] <= r_data[8499];
                
                r_data[8501] <= r_data[8500];
                
                r_data[8502] <= r_data[8501];
                
                r_data[8503] <= r_data[8502];
                
                r_data[8504] <= r_data[8503];
                
                r_data[8505] <= r_data[8504];
                
                r_data[8506] <= r_data[8505];
                
                r_data[8507] <= r_data[8506];
                
                r_data[8508] <= r_data[8507];
                
                r_data[8509] <= r_data[8508];
                
                r_data[8510] <= r_data[8509];
                
                r_data[8511] <= r_data[8510];
                
                r_data[8512] <= r_data[8511];
                
                r_data[8513] <= r_data[8512];
                
                r_data[8514] <= r_data[8513];
                
                r_data[8515] <= r_data[8514];
                
                r_data[8516] <= r_data[8515];
                
                r_data[8517] <= r_data[8516];
                
                r_data[8518] <= r_data[8517];
                
                r_data[8519] <= r_data[8518];
                
                r_data[8520] <= r_data[8519];
                
                r_data[8521] <= r_data[8520];
                
                r_data[8522] <= r_data[8521];
                
                r_data[8523] <= r_data[8522];
                
                r_data[8524] <= r_data[8523];
                
                r_data[8525] <= r_data[8524];
                
                r_data[8526] <= r_data[8525];
                
                r_data[8527] <= r_data[8526];
                
                r_data[8528] <= r_data[8527];
                
                r_data[8529] <= r_data[8528];
                
                r_data[8530] <= r_data[8529];
                
                r_data[8531] <= r_data[8530];
                
                r_data[8532] <= r_data[8531];
                
                r_data[8533] <= r_data[8532];
                
                r_data[8534] <= r_data[8533];
                
                r_data[8535] <= r_data[8534];
                
                r_data[8536] <= r_data[8535];
                
                r_data[8537] <= r_data[8536];
                
                r_data[8538] <= r_data[8537];
                
                r_data[8539] <= r_data[8538];
                
                r_data[8540] <= r_data[8539];
                
                r_data[8541] <= r_data[8540];
                
                r_data[8542] <= r_data[8541];
                
                r_data[8543] <= r_data[8542];
                
                r_data[8544] <= r_data[8543];
                
                r_data[8545] <= r_data[8544];
                
                r_data[8546] <= r_data[8545];
                
                r_data[8547] <= r_data[8546];
                
                r_data[8548] <= r_data[8547];
                
                r_data[8549] <= r_data[8548];
                
                r_data[8550] <= r_data[8549];
                
                r_data[8551] <= r_data[8550];
                
                r_data[8552] <= r_data[8551];
                
                r_data[8553] <= r_data[8552];
                
                r_data[8554] <= r_data[8553];
                
                r_data[8555] <= r_data[8554];
                
                r_data[8556] <= r_data[8555];
                
                r_data[8557] <= r_data[8556];
                
                r_data[8558] <= r_data[8557];
                
                r_data[8559] <= r_data[8558];
                
                r_data[8560] <= r_data[8559];
                
                r_data[8561] <= r_data[8560];
                
                r_data[8562] <= r_data[8561];
                
                r_data[8563] <= r_data[8562];
                
                r_data[8564] <= r_data[8563];
                
                r_data[8565] <= r_data[8564];
                
                r_data[8566] <= r_data[8565];
                
                r_data[8567] <= r_data[8566];
                
                r_data[8568] <= r_data[8567];
                
                r_data[8569] <= r_data[8568];
                
                r_data[8570] <= r_data[8569];
                
                r_data[8571] <= r_data[8570];
                
                r_data[8572] <= r_data[8571];
                
                r_data[8573] <= r_data[8572];
                
                r_data[8574] <= r_data[8573];
                
                r_data[8575] <= r_data[8574];
                
                r_data[8576] <= r_data[8575];
                
                r_data[8577] <= r_data[8576];
                
                r_data[8578] <= r_data[8577];
                
                r_data[8579] <= r_data[8578];
                
                r_data[8580] <= r_data[8579];
                
                r_data[8581] <= r_data[8580];
                
                r_data[8582] <= r_data[8581];
                
                r_data[8583] <= r_data[8582];
                
                r_data[8584] <= r_data[8583];
                
                r_data[8585] <= r_data[8584];
                
                r_data[8586] <= r_data[8585];
                
                r_data[8587] <= r_data[8586];
                
                r_data[8588] <= r_data[8587];
                
                r_data[8589] <= r_data[8588];
                
                r_data[8590] <= r_data[8589];
                
                r_data[8591] <= r_data[8590];
                
                r_data[8592] <= r_data[8591];
                
                r_data[8593] <= r_data[8592];
                
                r_data[8594] <= r_data[8593];
                
                r_data[8595] <= r_data[8594];
                
                r_data[8596] <= r_data[8595];
                
                r_data[8597] <= r_data[8596];
                
                r_data[8598] <= r_data[8597];
                
                r_data[8599] <= r_data[8598];
                
                r_data[8600] <= r_data[8599];
                
                r_data[8601] <= r_data[8600];
                
                r_data[8602] <= r_data[8601];
                
                r_data[8603] <= r_data[8602];
                
                r_data[8604] <= r_data[8603];
                
                r_data[8605] <= r_data[8604];
                
                r_data[8606] <= r_data[8605];
                
                r_data[8607] <= r_data[8606];
                
                r_data[8608] <= r_data[8607];
                
                r_data[8609] <= r_data[8608];
                
                r_data[8610] <= r_data[8609];
                
                r_data[8611] <= r_data[8610];
                
                r_data[8612] <= r_data[8611];
                
                r_data[8613] <= r_data[8612];
                
                r_data[8614] <= r_data[8613];
                
                r_data[8615] <= r_data[8614];
                
                r_data[8616] <= r_data[8615];
                
                r_data[8617] <= r_data[8616];
                
                r_data[8618] <= r_data[8617];
                
                r_data[8619] <= r_data[8618];
                
                r_data[8620] <= r_data[8619];
                
                r_data[8621] <= r_data[8620];
                
                r_data[8622] <= r_data[8621];
                
                r_data[8623] <= r_data[8622];
                
                r_data[8624] <= r_data[8623];
                
                r_data[8625] <= r_data[8624];
                
                r_data[8626] <= r_data[8625];
                
                r_data[8627] <= r_data[8626];
                
                r_data[8628] <= r_data[8627];
                
                r_data[8629] <= r_data[8628];
                
                r_data[8630] <= r_data[8629];
                
                r_data[8631] <= r_data[8630];
                
                r_data[8632] <= r_data[8631];
                
                r_data[8633] <= r_data[8632];
                
                r_data[8634] <= r_data[8633];
                
                r_data[8635] <= r_data[8634];
                
                r_data[8636] <= r_data[8635];
                
                r_data[8637] <= r_data[8636];
                
                r_data[8638] <= r_data[8637];
                
                r_data[8639] <= r_data[8638];
                
                r_data[8640] <= r_data[8639];
                
                r_data[8641] <= r_data[8640];
                
                r_data[8642] <= r_data[8641];
                
                r_data[8643] <= r_data[8642];
                
                r_data[8644] <= r_data[8643];
                
                r_data[8645] <= r_data[8644];
                
                r_data[8646] <= r_data[8645];
                
                r_data[8647] <= r_data[8646];
                
                r_data[8648] <= r_data[8647];
                
                r_data[8649] <= r_data[8648];
                
                r_data[8650] <= r_data[8649];
                
                r_data[8651] <= r_data[8650];
                
                r_data[8652] <= r_data[8651];
                
                r_data[8653] <= r_data[8652];
                
                r_data[8654] <= r_data[8653];
                
                r_data[8655] <= r_data[8654];
                
                r_data[8656] <= r_data[8655];
                
                r_data[8657] <= r_data[8656];
                
                r_data[8658] <= r_data[8657];
                
                r_data[8659] <= r_data[8658];
                
                r_data[8660] <= r_data[8659];
                
                r_data[8661] <= r_data[8660];
                
                r_data[8662] <= r_data[8661];
                
                r_data[8663] <= r_data[8662];
                
                r_data[8664] <= r_data[8663];
                
                r_data[8665] <= r_data[8664];
                
                r_data[8666] <= r_data[8665];
                
                r_data[8667] <= r_data[8666];
                
                r_data[8668] <= r_data[8667];
                
                r_data[8669] <= r_data[8668];
                
                r_data[8670] <= r_data[8669];
                
                r_data[8671] <= r_data[8670];
                
                r_data[8672] <= r_data[8671];
                
                r_data[8673] <= r_data[8672];
                
                r_data[8674] <= r_data[8673];
                
                r_data[8675] <= r_data[8674];
                
                r_data[8676] <= r_data[8675];
                
                r_data[8677] <= r_data[8676];
                
                r_data[8678] <= r_data[8677];
                
                r_data[8679] <= r_data[8678];
                
                r_data[8680] <= r_data[8679];
                
                r_data[8681] <= r_data[8680];
                
                r_data[8682] <= r_data[8681];
                
                r_data[8683] <= r_data[8682];
                
                r_data[8684] <= r_data[8683];
                
                r_data[8685] <= r_data[8684];
                
                r_data[8686] <= r_data[8685];
                
                r_data[8687] <= r_data[8686];
                
                r_data[8688] <= r_data[8687];
                
                r_data[8689] <= r_data[8688];
                
                r_data[8690] <= r_data[8689];
                
                r_data[8691] <= r_data[8690];
                
                r_data[8692] <= r_data[8691];
                
                r_data[8693] <= r_data[8692];
                
                r_data[8694] <= r_data[8693];
                
                r_data[8695] <= r_data[8694];
                
                r_data[8696] <= r_data[8695];
                
                r_data[8697] <= r_data[8696];
                
                r_data[8698] <= r_data[8697];
                
                r_data[8699] <= r_data[8698];
                
                r_data[8700] <= r_data[8699];
                
                r_data[8701] <= r_data[8700];
                
                r_data[8702] <= r_data[8701];
                
                r_data[8703] <= r_data[8702];
                
                r_data[8704] <= r_data[8703];
                
                r_data[8705] <= r_data[8704];
                
                r_data[8706] <= r_data[8705];
                
                r_data[8707] <= r_data[8706];
                
                r_data[8708] <= r_data[8707];
                
                r_data[8709] <= r_data[8708];
                
                r_data[8710] <= r_data[8709];
                
                r_data[8711] <= r_data[8710];
                
                r_data[8712] <= r_data[8711];
                
                r_data[8713] <= r_data[8712];
                
                r_data[8714] <= r_data[8713];
                
                r_data[8715] <= r_data[8714];
                
                r_data[8716] <= r_data[8715];
                
                r_data[8717] <= r_data[8716];
                
                r_data[8718] <= r_data[8717];
                
                r_data[8719] <= r_data[8718];
                
                r_data[8720] <= r_data[8719];
                
                r_data[8721] <= r_data[8720];
                
                r_data[8722] <= r_data[8721];
                
                r_data[8723] <= r_data[8722];
                
                r_data[8724] <= r_data[8723];
                
                r_data[8725] <= r_data[8724];
                
                r_data[8726] <= r_data[8725];
                
                r_data[8727] <= r_data[8726];
                
                r_data[8728] <= r_data[8727];
                
                r_data[8729] <= r_data[8728];
                
                r_data[8730] <= r_data[8729];
                
                r_data[8731] <= r_data[8730];
                
                r_data[8732] <= r_data[8731];
                
                r_data[8733] <= r_data[8732];
                
                r_data[8734] <= r_data[8733];
                
                r_data[8735] <= r_data[8734];
                
                r_data[8736] <= r_data[8735];
                
                r_data[8737] <= r_data[8736];
                
                r_data[8738] <= r_data[8737];
                
                r_data[8739] <= r_data[8738];
                
                r_data[8740] <= r_data[8739];
                
                r_data[8741] <= r_data[8740];
                
                r_data[8742] <= r_data[8741];
                
                r_data[8743] <= r_data[8742];
                
                r_data[8744] <= r_data[8743];
                
                r_data[8745] <= r_data[8744];
                
                r_data[8746] <= r_data[8745];
                
                r_data[8747] <= r_data[8746];
                
                r_data[8748] <= r_data[8747];
                
                r_data[8749] <= r_data[8748];
                
                r_data[8750] <= r_data[8749];
                
                r_data[8751] <= r_data[8750];
                
                r_data[8752] <= r_data[8751];
                
                r_data[8753] <= r_data[8752];
                
                r_data[8754] <= r_data[8753];
                
                r_data[8755] <= r_data[8754];
                
                r_data[8756] <= r_data[8755];
                
                r_data[8757] <= r_data[8756];
                
                r_data[8758] <= r_data[8757];
                
                r_data[8759] <= r_data[8758];
                
                r_data[8760] <= r_data[8759];
                
                r_data[8761] <= r_data[8760];
                
                r_data[8762] <= r_data[8761];
                
                r_data[8763] <= r_data[8762];
                
                r_data[8764] <= r_data[8763];
                
                r_data[8765] <= r_data[8764];
                
                r_data[8766] <= r_data[8765];
                
                r_data[8767] <= r_data[8766];
                
                r_data[8768] <= r_data[8767];
                
                r_data[8769] <= r_data[8768];
                
                r_data[8770] <= r_data[8769];
                
                r_data[8771] <= r_data[8770];
                
                r_data[8772] <= r_data[8771];
                
                r_data[8773] <= r_data[8772];
                
                r_data[8774] <= r_data[8773];
                
                r_data[8775] <= r_data[8774];
                
                r_data[8776] <= r_data[8775];
                
                r_data[8777] <= r_data[8776];
                
                r_data[8778] <= r_data[8777];
                
                r_data[8779] <= r_data[8778];
                
                r_data[8780] <= r_data[8779];
                
                r_data[8781] <= r_data[8780];
                
                r_data[8782] <= r_data[8781];
                
                r_data[8783] <= r_data[8782];
                
                r_data[8784] <= r_data[8783];
                
                r_data[8785] <= r_data[8784];
                
                r_data[8786] <= r_data[8785];
                
                r_data[8787] <= r_data[8786];
                
                r_data[8788] <= r_data[8787];
                
                r_data[8789] <= r_data[8788];
                
                r_data[8790] <= r_data[8789];
                
                r_data[8791] <= r_data[8790];
                
                r_data[8792] <= r_data[8791];
                
                r_data[8793] <= r_data[8792];
                
                r_data[8794] <= r_data[8793];
                
                r_data[8795] <= r_data[8794];
                
                r_data[8796] <= r_data[8795];
                
                r_data[8797] <= r_data[8796];
                
                r_data[8798] <= r_data[8797];
                
                r_data[8799] <= r_data[8798];
                
                r_data[8800] <= r_data[8799];
                
                r_data[8801] <= r_data[8800];
                
                r_data[8802] <= r_data[8801];
                
                r_data[8803] <= r_data[8802];
                
                r_data[8804] <= r_data[8803];
                
                r_data[8805] <= r_data[8804];
                
                r_data[8806] <= r_data[8805];
                
                r_data[8807] <= r_data[8806];
                
                r_data[8808] <= r_data[8807];
                
                r_data[8809] <= r_data[8808];
                
                r_data[8810] <= r_data[8809];
                
                r_data[8811] <= r_data[8810];
                
                r_data[8812] <= r_data[8811];
                
                r_data[8813] <= r_data[8812];
                
                r_data[8814] <= r_data[8813];
                
                r_data[8815] <= r_data[8814];
                
                r_data[8816] <= r_data[8815];
                
                r_data[8817] <= r_data[8816];
                
                r_data[8818] <= r_data[8817];
                
                r_data[8819] <= r_data[8818];
                
                r_data[8820] <= r_data[8819];
                
                r_data[8821] <= r_data[8820];
                
                r_data[8822] <= r_data[8821];
                
                r_data[8823] <= r_data[8822];
                
                r_data[8824] <= r_data[8823];
                
                r_data[8825] <= r_data[8824];
                
                r_data[8826] <= r_data[8825];
                
                r_data[8827] <= r_data[8826];
                
                r_data[8828] <= r_data[8827];
                
                r_data[8829] <= r_data[8828];
                
                r_data[8830] <= r_data[8829];
                
                r_data[8831] <= r_data[8830];
                
                r_data[8832] <= r_data[8831];
                
                r_data[8833] <= r_data[8832];
                
                r_data[8834] <= r_data[8833];
                
                r_data[8835] <= r_data[8834];
                
                r_data[8836] <= r_data[8835];
                
                r_data[8837] <= r_data[8836];
                
                r_data[8838] <= r_data[8837];
                
                r_data[8839] <= r_data[8838];
                
                r_data[8840] <= r_data[8839];
                
                r_data[8841] <= r_data[8840];
                
                r_data[8842] <= r_data[8841];
                
                r_data[8843] <= r_data[8842];
                
                r_data[8844] <= r_data[8843];
                
                r_data[8845] <= r_data[8844];
                
                r_data[8846] <= r_data[8845];
                
                r_data[8847] <= r_data[8846];
                
                r_data[8848] <= r_data[8847];
                
                r_data[8849] <= r_data[8848];
                
                r_data[8850] <= r_data[8849];
                
                r_data[8851] <= r_data[8850];
                
                r_data[8852] <= r_data[8851];
                
                r_data[8853] <= r_data[8852];
                
                r_data[8854] <= r_data[8853];
                
                r_data[8855] <= r_data[8854];
                
                r_data[8856] <= r_data[8855];
                
                r_data[8857] <= r_data[8856];
                
                r_data[8858] <= r_data[8857];
                
                r_data[8859] <= r_data[8858];
                
                r_data[8860] <= r_data[8859];
                
                r_data[8861] <= r_data[8860];
                
                r_data[8862] <= r_data[8861];
                
                r_data[8863] <= r_data[8862];
                
                r_data[8864] <= r_data[8863];
                
                r_data[8865] <= r_data[8864];
                
                r_data[8866] <= r_data[8865];
                
                r_data[8867] <= r_data[8866];
                
                r_data[8868] <= r_data[8867];
                
                r_data[8869] <= r_data[8868];
                
                r_data[8870] <= r_data[8869];
                
                r_data[8871] <= r_data[8870];
                
                r_data[8872] <= r_data[8871];
                
                r_data[8873] <= r_data[8872];
                
                r_data[8874] <= r_data[8873];
                
                r_data[8875] <= r_data[8874];
                
                r_data[8876] <= r_data[8875];
                
                r_data[8877] <= r_data[8876];
                
                r_data[8878] <= r_data[8877];
                
                r_data[8879] <= r_data[8878];
                
                r_data[8880] <= r_data[8879];
                
                r_data[8881] <= r_data[8880];
                
                r_data[8882] <= r_data[8881];
                
                r_data[8883] <= r_data[8882];
                
                r_data[8884] <= r_data[8883];
                
                r_data[8885] <= r_data[8884];
                
                r_data[8886] <= r_data[8885];
                
                r_data[8887] <= r_data[8886];
                
                r_data[8888] <= r_data[8887];
                
                r_data[8889] <= r_data[8888];
                
                r_data[8890] <= r_data[8889];
                
                r_data[8891] <= r_data[8890];
                
                r_data[8892] <= r_data[8891];
                
                r_data[8893] <= r_data[8892];
                
                r_data[8894] <= r_data[8893];
                
                r_data[8895] <= r_data[8894];
                
                r_data[8896] <= r_data[8895];
                
                r_data[8897] <= r_data[8896];
                
                r_data[8898] <= r_data[8897];
                
                r_data[8899] <= r_data[8898];
                
                r_data[8900] <= r_data[8899];
                
                r_data[8901] <= r_data[8900];
                
                r_data[8902] <= r_data[8901];
                
                r_data[8903] <= r_data[8902];
                
                r_data[8904] <= r_data[8903];
                
                r_data[8905] <= r_data[8904];
                
                r_data[8906] <= r_data[8905];
                
                r_data[8907] <= r_data[8906];
                
                r_data[8908] <= r_data[8907];
                
                r_data[8909] <= r_data[8908];
                
                r_data[8910] <= r_data[8909];
                
                r_data[8911] <= r_data[8910];
                
                r_data[8912] <= r_data[8911];
                
                r_data[8913] <= r_data[8912];
                
                r_data[8914] <= r_data[8913];
                
                r_data[8915] <= r_data[8914];
                
                r_data[8916] <= r_data[8915];
                
                r_data[8917] <= r_data[8916];
                
                r_data[8918] <= r_data[8917];
                
                r_data[8919] <= r_data[8918];
                
                r_data[8920] <= r_data[8919];
                
                r_data[8921] <= r_data[8920];
                
                r_data[8922] <= r_data[8921];
                
                r_data[8923] <= r_data[8922];
                
                r_data[8924] <= r_data[8923];
                
                r_data[8925] <= r_data[8924];
                
                r_data[8926] <= r_data[8925];
                
                r_data[8927] <= r_data[8926];
                
                r_data[8928] <= r_data[8927];
                
                r_data[8929] <= r_data[8928];
                
                r_data[8930] <= r_data[8929];
                
                r_data[8931] <= r_data[8930];
                
                r_data[8932] <= r_data[8931];
                
                r_data[8933] <= r_data[8932];
                
                r_data[8934] <= r_data[8933];
                
                r_data[8935] <= r_data[8934];
                
                r_data[8936] <= r_data[8935];
                
                r_data[8937] <= r_data[8936];
                
                r_data[8938] <= r_data[8937];
                
                r_data[8939] <= r_data[8938];
                
                r_data[8940] <= r_data[8939];
                
                r_data[8941] <= r_data[8940];
                
                r_data[8942] <= r_data[8941];
                
                r_data[8943] <= r_data[8942];
                
                r_data[8944] <= r_data[8943];
                
                r_data[8945] <= r_data[8944];
                
                r_data[8946] <= r_data[8945];
                
                r_data[8947] <= r_data[8946];
                
                r_data[8948] <= r_data[8947];
                
                r_data[8949] <= r_data[8948];
                
                r_data[8950] <= r_data[8949];
                
                r_data[8951] <= r_data[8950];
                
                r_data[8952] <= r_data[8951];
                
                r_data[8953] <= r_data[8952];
                
                r_data[8954] <= r_data[8953];
                
                r_data[8955] <= r_data[8954];
                
                r_data[8956] <= r_data[8955];
                
                r_data[8957] <= r_data[8956];
                
                r_data[8958] <= r_data[8957];
                
                r_data[8959] <= r_data[8958];
                
                r_data[8960] <= r_data[8959];
                
                r_data[8961] <= r_data[8960];
                
                r_data[8962] <= r_data[8961];
                
                r_data[8963] <= r_data[8962];
                
                r_data[8964] <= r_data[8963];
                
                r_data[8965] <= r_data[8964];
                
                r_data[8966] <= r_data[8965];
                
                r_data[8967] <= r_data[8966];
                
                r_data[8968] <= r_data[8967];
                
                r_data[8969] <= r_data[8968];
                
                r_data[8970] <= r_data[8969];
                
                r_data[8971] <= r_data[8970];
                
                r_data[8972] <= r_data[8971];
                
                r_data[8973] <= r_data[8972];
                
                r_data[8974] <= r_data[8973];
                
                r_data[8975] <= r_data[8974];
                
                r_data[8976] <= r_data[8975];
                
                r_data[8977] <= r_data[8976];
                
                r_data[8978] <= r_data[8977];
                
                r_data[8979] <= r_data[8978];
                
                r_data[8980] <= r_data[8979];
                
                r_data[8981] <= r_data[8980];
                
                r_data[8982] <= r_data[8981];
                
                r_data[8983] <= r_data[8982];
                
                r_data[8984] <= r_data[8983];
                
                r_data[8985] <= r_data[8984];
                
                r_data[8986] <= r_data[8985];
                
                r_data[8987] <= r_data[8986];
                
                r_data[8988] <= r_data[8987];
                
                r_data[8989] <= r_data[8988];
                
                r_data[8990] <= r_data[8989];
                
                r_data[8991] <= r_data[8990];
                
                r_data[8992] <= r_data[8991];
                
                r_data[8993] <= r_data[8992];
                
                r_data[8994] <= r_data[8993];
                
                r_data[8995] <= r_data[8994];
                
                r_data[8996] <= r_data[8995];
                
                r_data[8997] <= r_data[8996];
                
                r_data[8998] <= r_data[8997];
                
                r_data[8999] <= r_data[8998];
                
                r_data[9000] <= r_data[8999];
                
                r_data[9001] <= r_data[9000];
                
                r_data[9002] <= r_data[9001];
                
                r_data[9003] <= r_data[9002];
                
                r_data[9004] <= r_data[9003];
                
                r_data[9005] <= r_data[9004];
                
                r_data[9006] <= r_data[9005];
                
                r_data[9007] <= r_data[9006];
                
                r_data[9008] <= r_data[9007];
                
                r_data[9009] <= r_data[9008];
                
                r_data[9010] <= r_data[9009];
                
                r_data[9011] <= r_data[9010];
                
                r_data[9012] <= r_data[9011];
                
                r_data[9013] <= r_data[9012];
                
                r_data[9014] <= r_data[9013];
                
                r_data[9015] <= r_data[9014];
                
                r_data[9016] <= r_data[9015];
                
                r_data[9017] <= r_data[9016];
                
                r_data[9018] <= r_data[9017];
                
                r_data[9019] <= r_data[9018];
                
                r_data[9020] <= r_data[9019];
                
                r_data[9021] <= r_data[9020];
                
                r_data[9022] <= r_data[9021];
                
                r_data[9023] <= r_data[9022];
                
                r_data[9024] <= r_data[9023];
                
                r_data[9025] <= r_data[9024];
                
                r_data[9026] <= r_data[9025];
                
                r_data[9027] <= r_data[9026];
                
                r_data[9028] <= r_data[9027];
                
                r_data[9029] <= r_data[9028];
                
                r_data[9030] <= r_data[9029];
                
                r_data[9031] <= r_data[9030];
                
                r_data[9032] <= r_data[9031];
                
                r_data[9033] <= r_data[9032];
                
                r_data[9034] <= r_data[9033];
                
                r_data[9035] <= r_data[9034];
                
                r_data[9036] <= r_data[9035];
                
                r_data[9037] <= r_data[9036];
                
                r_data[9038] <= r_data[9037];
                
                r_data[9039] <= r_data[9038];
                
                r_data[9040] <= r_data[9039];
                
                r_data[9041] <= r_data[9040];
                
                r_data[9042] <= r_data[9041];
                
                r_data[9043] <= r_data[9042];
                
                r_data[9044] <= r_data[9043];
                
                r_data[9045] <= r_data[9044];
                
                r_data[9046] <= r_data[9045];
                
                r_data[9047] <= r_data[9046];
                
                r_data[9048] <= r_data[9047];
                
                r_data[9049] <= r_data[9048];
                
                r_data[9050] <= r_data[9049];
                
                r_data[9051] <= r_data[9050];
                
                r_data[9052] <= r_data[9051];
                
                r_data[9053] <= r_data[9052];
                
                r_data[9054] <= r_data[9053];
                
                r_data[9055] <= r_data[9054];
                
                r_data[9056] <= r_data[9055];
                
                r_data[9057] <= r_data[9056];
                
                r_data[9058] <= r_data[9057];
                
                r_data[9059] <= r_data[9058];
                
                r_data[9060] <= r_data[9059];
                
                r_data[9061] <= r_data[9060];
                
                r_data[9062] <= r_data[9061];
                
                r_data[9063] <= r_data[9062];
                
                r_data[9064] <= r_data[9063];
                
                r_data[9065] <= r_data[9064];
                
                r_data[9066] <= r_data[9065];
                
                r_data[9067] <= r_data[9066];
                
                r_data[9068] <= r_data[9067];
                
                r_data[9069] <= r_data[9068];
                
                r_data[9070] <= r_data[9069];
                
                r_data[9071] <= r_data[9070];
                
                r_data[9072] <= r_data[9071];
                
                r_data[9073] <= r_data[9072];
                
                r_data[9074] <= r_data[9073];
                
                r_data[9075] <= r_data[9074];
                
                r_data[9076] <= r_data[9075];
                
                r_data[9077] <= r_data[9076];
                
                r_data[9078] <= r_data[9077];
                
                r_data[9079] <= r_data[9078];
                
                r_data[9080] <= r_data[9079];
                
                r_data[9081] <= r_data[9080];
                
                r_data[9082] <= r_data[9081];
                
                r_data[9083] <= r_data[9082];
                
                r_data[9084] <= r_data[9083];
                
                r_data[9085] <= r_data[9084];
                
                r_data[9086] <= r_data[9085];
                
                r_data[9087] <= r_data[9086];
                
                r_data[9088] <= r_data[9087];
                
                r_data[9089] <= r_data[9088];
                
                r_data[9090] <= r_data[9089];
                
                r_data[9091] <= r_data[9090];
                
                r_data[9092] <= r_data[9091];
                
                r_data[9093] <= r_data[9092];
                
                r_data[9094] <= r_data[9093];
                
                r_data[9095] <= r_data[9094];
                
                r_data[9096] <= r_data[9095];
                
                r_data[9097] <= r_data[9096];
                
                r_data[9098] <= r_data[9097];
                
                r_data[9099] <= r_data[9098];
                
                r_data[9100] <= r_data[9099];
                
                r_data[9101] <= r_data[9100];
                
                r_data[9102] <= r_data[9101];
                
                r_data[9103] <= r_data[9102];
                
                r_data[9104] <= r_data[9103];
                
                r_data[9105] <= r_data[9104];
                
                r_data[9106] <= r_data[9105];
                
                r_data[9107] <= r_data[9106];
                
                r_data[9108] <= r_data[9107];
                
                r_data[9109] <= r_data[9108];
                
                r_data[9110] <= r_data[9109];
                
                r_data[9111] <= r_data[9110];
                
                r_data[9112] <= r_data[9111];
                
                r_data[9113] <= r_data[9112];
                
                r_data[9114] <= r_data[9113];
                
                r_data[9115] <= r_data[9114];
                
                r_data[9116] <= r_data[9115];
                
                r_data[9117] <= r_data[9116];
                
                r_data[9118] <= r_data[9117];
                
                r_data[9119] <= r_data[9118];
                
                r_data[9120] <= r_data[9119];
                
                r_data[9121] <= r_data[9120];
                
                r_data[9122] <= r_data[9121];
                
                r_data[9123] <= r_data[9122];
                
                r_data[9124] <= r_data[9123];
                
                r_data[9125] <= r_data[9124];
                
                r_data[9126] <= r_data[9125];
                
                r_data[9127] <= r_data[9126];
                
                r_data[9128] <= r_data[9127];
                
                r_data[9129] <= r_data[9128];
                
                r_data[9130] <= r_data[9129];
                
                r_data[9131] <= r_data[9130];
                
                r_data[9132] <= r_data[9131];
                
                r_data[9133] <= r_data[9132];
                
                r_data[9134] <= r_data[9133];
                
                r_data[9135] <= r_data[9134];
                
                r_data[9136] <= r_data[9135];
                
                r_data[9137] <= r_data[9136];
                
                r_data[9138] <= r_data[9137];
                
                r_data[9139] <= r_data[9138];
                
                r_data[9140] <= r_data[9139];
                
                r_data[9141] <= r_data[9140];
                
                r_data[9142] <= r_data[9141];
                
                r_data[9143] <= r_data[9142];
                
                r_data[9144] <= r_data[9143];
                
                r_data[9145] <= r_data[9144];
                
                r_data[9146] <= r_data[9145];
                
                r_data[9147] <= r_data[9146];
                
                r_data[9148] <= r_data[9147];
                
                r_data[9149] <= r_data[9148];
                
                r_data[9150] <= r_data[9149];
                
                r_data[9151] <= r_data[9150];
                
                r_data[9152] <= r_data[9151];
                
                r_data[9153] <= r_data[9152];
                
                r_data[9154] <= r_data[9153];
                
                r_data[9155] <= r_data[9154];
                
                r_data[9156] <= r_data[9155];
                
                r_data[9157] <= r_data[9156];
                
                r_data[9158] <= r_data[9157];
                
                r_data[9159] <= r_data[9158];
                
                r_data[9160] <= r_data[9159];
                
                r_data[9161] <= r_data[9160];
                
                r_data[9162] <= r_data[9161];
                
                r_data[9163] <= r_data[9162];
                
                r_data[9164] <= r_data[9163];
                
                r_data[9165] <= r_data[9164];
                
                r_data[9166] <= r_data[9165];
                
                r_data[9167] <= r_data[9166];
                
                r_data[9168] <= r_data[9167];
                
                r_data[9169] <= r_data[9168];
                
                r_data[9170] <= r_data[9169];
                
                r_data[9171] <= r_data[9170];
                
                r_data[9172] <= r_data[9171];
                
                r_data[9173] <= r_data[9172];
                
                r_data[9174] <= r_data[9173];
                
                r_data[9175] <= r_data[9174];
                
                r_data[9176] <= r_data[9175];
                
                r_data[9177] <= r_data[9176];
                
                r_data[9178] <= r_data[9177];
                
                r_data[9179] <= r_data[9178];
                
                r_data[9180] <= r_data[9179];
                
                r_data[9181] <= r_data[9180];
                
                r_data[9182] <= r_data[9181];
                
                r_data[9183] <= r_data[9182];
                
                r_data[9184] <= r_data[9183];
                
                r_data[9185] <= r_data[9184];
                
                r_data[9186] <= r_data[9185];
                
                r_data[9187] <= r_data[9186];
                
                r_data[9188] <= r_data[9187];
                
                r_data[9189] <= r_data[9188];
                
                r_data[9190] <= r_data[9189];
                
                r_data[9191] <= r_data[9190];
                
                r_data[9192] <= r_data[9191];
                
                r_data[9193] <= r_data[9192];
                
                r_data[9194] <= r_data[9193];
                
                r_data[9195] <= r_data[9194];
                
                r_data[9196] <= r_data[9195];
                
                r_data[9197] <= r_data[9196];
                
                r_data[9198] <= r_data[9197];
                
                r_data[9199] <= r_data[9198];
                
                r_data[9200] <= r_data[9199];
                
                r_data[9201] <= r_data[9200];
                
                r_data[9202] <= r_data[9201];
                
                r_data[9203] <= r_data[9202];
                
                r_data[9204] <= r_data[9203];
                
                r_data[9205] <= r_data[9204];
                
                r_data[9206] <= r_data[9205];
                
                r_data[9207] <= r_data[9206];
                
                r_data[9208] <= r_data[9207];
                
                r_data[9209] <= r_data[9208];
                
                r_data[9210] <= r_data[9209];
                
                r_data[9211] <= r_data[9210];
                
                r_data[9212] <= r_data[9211];
                
                r_data[9213] <= r_data[9212];
                
                r_data[9214] <= r_data[9213];
                
                r_data[9215] <= r_data[9214];
                
                r_data[9216] <= r_data[9215];
                
                r_data[9217] <= r_data[9216];
                
                r_data[9218] <= r_data[9217];
                
                r_data[9219] <= r_data[9218];
                
                r_data[9220] <= r_data[9219];
                
                r_data[9221] <= r_data[9220];
                
                r_data[9222] <= r_data[9221];
                
                r_data[9223] <= r_data[9222];
                
                r_data[9224] <= r_data[9223];
                
                r_data[9225] <= r_data[9224];
                
                r_data[9226] <= r_data[9225];
                
                r_data[9227] <= r_data[9226];
                
                r_data[9228] <= r_data[9227];
                
                r_data[9229] <= r_data[9228];
                
                r_data[9230] <= r_data[9229];
                
                r_data[9231] <= r_data[9230];
                
                r_data[9232] <= r_data[9231];
                
                r_data[9233] <= r_data[9232];
                
                r_data[9234] <= r_data[9233];
                
                r_data[9235] <= r_data[9234];
                
                r_data[9236] <= r_data[9235];
                
                r_data[9237] <= r_data[9236];
                
                r_data[9238] <= r_data[9237];
                
                r_data[9239] <= r_data[9238];
                
                r_data[9240] <= r_data[9239];
                
                r_data[9241] <= r_data[9240];
                
                r_data[9242] <= r_data[9241];
                
                r_data[9243] <= r_data[9242];
                
                r_data[9244] <= r_data[9243];
                
                r_data[9245] <= r_data[9244];
                
                r_data[9246] <= r_data[9245];
                
                r_data[9247] <= r_data[9246];
                
                r_data[9248] <= r_data[9247];
                
                r_data[9249] <= r_data[9248];
                
                r_data[9250] <= r_data[9249];
                
                r_data[9251] <= r_data[9250];
                
                r_data[9252] <= r_data[9251];
                
                r_data[9253] <= r_data[9252];
                
                r_data[9254] <= r_data[9253];
                
                r_data[9255] <= r_data[9254];
                
                r_data[9256] <= r_data[9255];
                
                r_data[9257] <= r_data[9256];
                
                r_data[9258] <= r_data[9257];
                
                r_data[9259] <= r_data[9258];
                
                r_data[9260] <= r_data[9259];
                
                r_data[9261] <= r_data[9260];
                
                r_data[9262] <= r_data[9261];
                
                r_data[9263] <= r_data[9262];
                
                r_data[9264] <= r_data[9263];
                
                r_data[9265] <= r_data[9264];
                
                r_data[9266] <= r_data[9265];
                
                r_data[9267] <= r_data[9266];
                
                r_data[9268] <= r_data[9267];
                
                r_data[9269] <= r_data[9268];
                
                r_data[9270] <= r_data[9269];
                
                r_data[9271] <= r_data[9270];
                
                r_data[9272] <= r_data[9271];
                
                r_data[9273] <= r_data[9272];
                
                r_data[9274] <= r_data[9273];
                
                r_data[9275] <= r_data[9274];
                
                r_data[9276] <= r_data[9275];
                
                r_data[9277] <= r_data[9276];
                
                r_data[9278] <= r_data[9277];
                
                r_data[9279] <= r_data[9278];
                
                r_data[9280] <= r_data[9279];
                
                r_data[9281] <= r_data[9280];
                
                r_data[9282] <= r_data[9281];
                
                r_data[9283] <= r_data[9282];
                
                r_data[9284] <= r_data[9283];
                
                r_data[9285] <= r_data[9284];
                
                r_data[9286] <= r_data[9285];
                
                r_data[9287] <= r_data[9286];
                
                r_data[9288] <= r_data[9287];
                
                r_data[9289] <= r_data[9288];
                
                r_data[9290] <= r_data[9289];
                
                r_data[9291] <= r_data[9290];
                
                r_data[9292] <= r_data[9291];
                
                r_data[9293] <= r_data[9292];
                
                r_data[9294] <= r_data[9293];
                
                r_data[9295] <= r_data[9294];
                
                r_data[9296] <= r_data[9295];
                
                r_data[9297] <= r_data[9296];
                
                r_data[9298] <= r_data[9297];
                
                r_data[9299] <= r_data[9298];
                
                r_data[9300] <= r_data[9299];
                
                r_data[9301] <= r_data[9300];
                
                r_data[9302] <= r_data[9301];
                
                r_data[9303] <= r_data[9302];
                
                r_data[9304] <= r_data[9303];
                
                r_data[9305] <= r_data[9304];
                
                r_data[9306] <= r_data[9305];
                
                r_data[9307] <= r_data[9306];
                
                r_data[9308] <= r_data[9307];
                
                r_data[9309] <= r_data[9308];
                
                r_data[9310] <= r_data[9309];
                
                r_data[9311] <= r_data[9310];
                
                r_data[9312] <= r_data[9311];
                
                r_data[9313] <= r_data[9312];
                
                r_data[9314] <= r_data[9313];
                
                r_data[9315] <= r_data[9314];
                
                r_data[9316] <= r_data[9315];
                
                r_data[9317] <= r_data[9316];
                
                r_data[9318] <= r_data[9317];
                
                r_data[9319] <= r_data[9318];
                
                r_data[9320] <= r_data[9319];
                
                r_data[9321] <= r_data[9320];
                
                r_data[9322] <= r_data[9321];
                
                r_data[9323] <= r_data[9322];
                
                r_data[9324] <= r_data[9323];
                
                r_data[9325] <= r_data[9324];
                
                r_data[9326] <= r_data[9325];
                
                r_data[9327] <= r_data[9326];
                
                r_data[9328] <= r_data[9327];
                
                r_data[9329] <= r_data[9328];
                
                r_data[9330] <= r_data[9329];
                
                r_data[9331] <= r_data[9330];
                
                r_data[9332] <= r_data[9331];
                
                r_data[9333] <= r_data[9332];
                
                r_data[9334] <= r_data[9333];
                
                r_data[9335] <= r_data[9334];
                
                r_data[9336] <= r_data[9335];
                
                r_data[9337] <= r_data[9336];
                
                r_data[9338] <= r_data[9337];
                
                r_data[9339] <= r_data[9338];
                
                r_data[9340] <= r_data[9339];
                
                r_data[9341] <= r_data[9340];
                
                r_data[9342] <= r_data[9341];
                
                r_data[9343] <= r_data[9342];
                
                r_data[9344] <= r_data[9343];
                
                r_data[9345] <= r_data[9344];
                
                r_data[9346] <= r_data[9345];
                
                r_data[9347] <= r_data[9346];
                
                r_data[9348] <= r_data[9347];
                
                r_data[9349] <= r_data[9348];
                
                r_data[9350] <= r_data[9349];
                
                r_data[9351] <= r_data[9350];
                
                r_data[9352] <= r_data[9351];
                
                r_data[9353] <= r_data[9352];
                
                r_data[9354] <= r_data[9353];
                
                r_data[9355] <= r_data[9354];
                
                r_data[9356] <= r_data[9355];
                
                r_data[9357] <= r_data[9356];
                
                r_data[9358] <= r_data[9357];
                
                r_data[9359] <= r_data[9358];
                
                r_data[9360] <= r_data[9359];
                
                r_data[9361] <= r_data[9360];
                
                r_data[9362] <= r_data[9361];
                
                r_data[9363] <= r_data[9362];
                
                r_data[9364] <= r_data[9363];
                
                r_data[9365] <= r_data[9364];
                
                r_data[9366] <= r_data[9365];
                
                r_data[9367] <= r_data[9366];
                
                r_data[9368] <= r_data[9367];
                
                r_data[9369] <= r_data[9368];
                
                r_data[9370] <= r_data[9369];
                
                r_data[9371] <= r_data[9370];
                
                r_data[9372] <= r_data[9371];
                
                r_data[9373] <= r_data[9372];
                
                r_data[9374] <= r_data[9373];
                
                r_data[9375] <= r_data[9374];
                
                r_data[9376] <= r_data[9375];
                
                r_data[9377] <= r_data[9376];
                
                r_data[9378] <= r_data[9377];
                
                r_data[9379] <= r_data[9378];
                
                r_data[9380] <= r_data[9379];
                
                r_data[9381] <= r_data[9380];
                
                r_data[9382] <= r_data[9381];
                
                r_data[9383] <= r_data[9382];
                
                r_data[9384] <= r_data[9383];
                
                r_data[9385] <= r_data[9384];
                
                r_data[9386] <= r_data[9385];
                
                r_data[9387] <= r_data[9386];
                
                r_data[9388] <= r_data[9387];
                
                r_data[9389] <= r_data[9388];
                
                r_data[9390] <= r_data[9389];
                
                r_data[9391] <= r_data[9390];
                
                r_data[9392] <= r_data[9391];
                
                r_data[9393] <= r_data[9392];
                
                r_data[9394] <= r_data[9393];
                
                r_data[9395] <= r_data[9394];
                
                r_data[9396] <= r_data[9395];
                
                r_data[9397] <= r_data[9396];
                
                r_data[9398] <= r_data[9397];
                
                r_data[9399] <= r_data[9398];
                
                r_data[9400] <= r_data[9399];
                
                r_data[9401] <= r_data[9400];
                
                r_data[9402] <= r_data[9401];
                
                r_data[9403] <= r_data[9402];
                
                r_data[9404] <= r_data[9403];
                
                r_data[9405] <= r_data[9404];
                
                r_data[9406] <= r_data[9405];
                
                r_data[9407] <= r_data[9406];
                
                r_data[9408] <= r_data[9407];
                
                r_data[9409] <= r_data[9408];
                
                r_data[9410] <= r_data[9409];
                
                r_data[9411] <= r_data[9410];
                
                r_data[9412] <= r_data[9411];
                
                r_data[9413] <= r_data[9412];
                
                r_data[9414] <= r_data[9413];
                
                r_data[9415] <= r_data[9414];
                
                r_data[9416] <= r_data[9415];
                
                r_data[9417] <= r_data[9416];
                
                r_data[9418] <= r_data[9417];
                
                r_data[9419] <= r_data[9418];
                
                r_data[9420] <= r_data[9419];
                
                r_data[9421] <= r_data[9420];
                
                r_data[9422] <= r_data[9421];
                
                r_data[9423] <= r_data[9422];
                
                r_data[9424] <= r_data[9423];
                
                r_data[9425] <= r_data[9424];
                
                r_data[9426] <= r_data[9425];
                
                r_data[9427] <= r_data[9426];
                
                r_data[9428] <= r_data[9427];
                
                r_data[9429] <= r_data[9428];
                
                r_data[9430] <= r_data[9429];
                
                r_data[9431] <= r_data[9430];
                
                r_data[9432] <= r_data[9431];
                
                r_data[9433] <= r_data[9432];
                
                r_data[9434] <= r_data[9433];
                
                r_data[9435] <= r_data[9434];
                
                r_data[9436] <= r_data[9435];
                
                r_data[9437] <= r_data[9436];
                
                r_data[9438] <= r_data[9437];
                
                r_data[9439] <= r_data[9438];
                
                r_data[9440] <= r_data[9439];
                
                r_data[9441] <= r_data[9440];
                
                r_data[9442] <= r_data[9441];
                
                r_data[9443] <= r_data[9442];
                
                r_data[9444] <= r_data[9443];
                
                r_data[9445] <= r_data[9444];
                
                r_data[9446] <= r_data[9445];
                
                r_data[9447] <= r_data[9446];
                
                r_data[9448] <= r_data[9447];
                
                r_data[9449] <= r_data[9448];
                
                r_data[9450] <= r_data[9449];
                
                r_data[9451] <= r_data[9450];
                
                r_data[9452] <= r_data[9451];
                
                r_data[9453] <= r_data[9452];
                
                r_data[9454] <= r_data[9453];
                
                r_data[9455] <= r_data[9454];
                
                r_data[9456] <= r_data[9455];
                
                r_data[9457] <= r_data[9456];
                
                r_data[9458] <= r_data[9457];
                
                r_data[9459] <= r_data[9458];
                
                r_data[9460] <= r_data[9459];
                
                r_data[9461] <= r_data[9460];
                
                r_data[9462] <= r_data[9461];
                
                r_data[9463] <= r_data[9462];
                
                r_data[9464] <= r_data[9463];
                
                r_data[9465] <= r_data[9464];
                
                r_data[9466] <= r_data[9465];
                
                r_data[9467] <= r_data[9466];
                
                r_data[9468] <= r_data[9467];
                
                r_data[9469] <= r_data[9468];
                
                r_data[9470] <= r_data[9469];
                
                r_data[9471] <= r_data[9470];
                
                r_data[9472] <= r_data[9471];
                
                r_data[9473] <= r_data[9472];
                
                r_data[9474] <= r_data[9473];
                
                r_data[9475] <= r_data[9474];
                
                r_data[9476] <= r_data[9475];
                
                r_data[9477] <= r_data[9476];
                
                r_data[9478] <= r_data[9477];
                
                r_data[9479] <= r_data[9478];
                
                r_data[9480] <= r_data[9479];
                
                r_data[9481] <= r_data[9480];
                
                r_data[9482] <= r_data[9481];
                
                r_data[9483] <= r_data[9482];
                
                r_data[9484] <= r_data[9483];
                
                r_data[9485] <= r_data[9484];
                
                r_data[9486] <= r_data[9485];
                
                r_data[9487] <= r_data[9486];
                
                r_data[9488] <= r_data[9487];
                
                r_data[9489] <= r_data[9488];
                
                r_data[9490] <= r_data[9489];
                
                r_data[9491] <= r_data[9490];
                
                r_data[9492] <= r_data[9491];
                
                r_data[9493] <= r_data[9492];
                
                r_data[9494] <= r_data[9493];
                
                r_data[9495] <= r_data[9494];
                
                r_data[9496] <= r_data[9495];
                
                r_data[9497] <= r_data[9496];
                
                r_data[9498] <= r_data[9497];
                
                r_data[9499] <= r_data[9498];
                
                r_data[9500] <= r_data[9499];
                
                r_data[9501] <= r_data[9500];
                
                r_data[9502] <= r_data[9501];
                
                r_data[9503] <= r_data[9502];
                
                r_data[9504] <= r_data[9503];
                
                r_data[9505] <= r_data[9504];
                
                r_data[9506] <= r_data[9505];
                
                r_data[9507] <= r_data[9506];
                
                r_data[9508] <= r_data[9507];
                
                r_data[9509] <= r_data[9508];
                
                r_data[9510] <= r_data[9509];
                
                r_data[9511] <= r_data[9510];
                
                r_data[9512] <= r_data[9511];
                
                r_data[9513] <= r_data[9512];
                
                r_data[9514] <= r_data[9513];
                
                r_data[9515] <= r_data[9514];
                
                r_data[9516] <= r_data[9515];
                
                r_data[9517] <= r_data[9516];
                
                r_data[9518] <= r_data[9517];
                
                r_data[9519] <= r_data[9518];
                
                r_data[9520] <= r_data[9519];
                
                r_data[9521] <= r_data[9520];
                
                r_data[9522] <= r_data[9521];
                
                r_data[9523] <= r_data[9522];
                
                r_data[9524] <= r_data[9523];
                
                r_data[9525] <= r_data[9524];
                
                r_data[9526] <= r_data[9525];
                
                r_data[9527] <= r_data[9526];
                
                r_data[9528] <= r_data[9527];
                
                r_data[9529] <= r_data[9528];
                
                r_data[9530] <= r_data[9529];
                
                r_data[9531] <= r_data[9530];
                
                r_data[9532] <= r_data[9531];
                
                r_data[9533] <= r_data[9532];
                
                r_data[9534] <= r_data[9533];
                
                r_data[9535] <= r_data[9534];
                
                r_data[9536] <= r_data[9535];
                
                r_data[9537] <= r_data[9536];
                
                r_data[9538] <= r_data[9537];
                
                r_data[9539] <= r_data[9538];
                
                r_data[9540] <= r_data[9539];
                
                r_data[9541] <= r_data[9540];
                
                r_data[9542] <= r_data[9541];
                
                r_data[9543] <= r_data[9542];
                
                r_data[9544] <= r_data[9543];
                
                r_data[9545] <= r_data[9544];
                
                r_data[9546] <= r_data[9545];
                
                r_data[9547] <= r_data[9546];
                
                r_data[9548] <= r_data[9547];
                
                r_data[9549] <= r_data[9548];
                
                r_data[9550] <= r_data[9549];
                
                r_data[9551] <= r_data[9550];
                
                r_data[9552] <= r_data[9551];
                
                r_data[9553] <= r_data[9552];
                
                r_data[9554] <= r_data[9553];
                
                r_data[9555] <= r_data[9554];
                
                r_data[9556] <= r_data[9555];
                
                r_data[9557] <= r_data[9556];
                
                r_data[9558] <= r_data[9557];
                
                r_data[9559] <= r_data[9558];
                
                r_data[9560] <= r_data[9559];
                
                r_data[9561] <= r_data[9560];
                
                r_data[9562] <= r_data[9561];
                
                r_data[9563] <= r_data[9562];
                
                r_data[9564] <= r_data[9563];
                
                r_data[9565] <= r_data[9564];
                
                r_data[9566] <= r_data[9565];
                
                r_data[9567] <= r_data[9566];
                
                r_data[9568] <= r_data[9567];
                
                r_data[9569] <= r_data[9568];
                
                r_data[9570] <= r_data[9569];
                
                r_data[9571] <= r_data[9570];
                
                r_data[9572] <= r_data[9571];
                
                r_data[9573] <= r_data[9572];
                
                r_data[9574] <= r_data[9573];
                
                r_data[9575] <= r_data[9574];
                
                r_data[9576] <= r_data[9575];
                
                r_data[9577] <= r_data[9576];
                
                r_data[9578] <= r_data[9577];
                
                r_data[9579] <= r_data[9578];
                
                r_data[9580] <= r_data[9579];
                
                r_data[9581] <= r_data[9580];
                
                r_data[9582] <= r_data[9581];
                
                r_data[9583] <= r_data[9582];
                
                r_data[9584] <= r_data[9583];
                
                r_data[9585] <= r_data[9584];
                
                r_data[9586] <= r_data[9585];
                
                r_data[9587] <= r_data[9586];
                
                r_data[9588] <= r_data[9587];
                
                r_data[9589] <= r_data[9588];
                
                r_data[9590] <= r_data[9589];
                
                r_data[9591] <= r_data[9590];
                
                r_data[9592] <= r_data[9591];
                
                r_data[9593] <= r_data[9592];
                
                r_data[9594] <= r_data[9593];
                
                r_data[9595] <= r_data[9594];
                
                r_data[9596] <= r_data[9595];
                
                r_data[9597] <= r_data[9596];
                
                r_data[9598] <= r_data[9597];
                
                r_data[9599] <= r_data[9598];
                
                r_data[9600] <= r_data[9599];
                
                r_data[9601] <= r_data[9600];
                
                r_data[9602] <= r_data[9601];
                
                r_data[9603] <= r_data[9602];
                
                r_data[9604] <= r_data[9603];
                
                r_data[9605] <= r_data[9604];
                
                r_data[9606] <= r_data[9605];
                
                r_data[9607] <= r_data[9606];
                
                r_data[9608] <= r_data[9607];
                
                r_data[9609] <= r_data[9608];
                
                r_data[9610] <= r_data[9609];
                
                r_data[9611] <= r_data[9610];
                
                r_data[9612] <= r_data[9611];
                
                r_data[9613] <= r_data[9612];
                
                r_data[9614] <= r_data[9613];
                
                r_data[9615] <= r_data[9614];
                
                r_data[9616] <= r_data[9615];
                
                r_data[9617] <= r_data[9616];
                
                r_data[9618] <= r_data[9617];
                
                r_data[9619] <= r_data[9618];
                
                r_data[9620] <= r_data[9619];
                
                r_data[9621] <= r_data[9620];
                
                r_data[9622] <= r_data[9621];
                
                r_data[9623] <= r_data[9622];
                
                r_data[9624] <= r_data[9623];
                
                r_data[9625] <= r_data[9624];
                
                r_data[9626] <= r_data[9625];
                
                r_data[9627] <= r_data[9626];
                
                r_data[9628] <= r_data[9627];
                
                r_data[9629] <= r_data[9628];
                
                r_data[9630] <= r_data[9629];
                
                r_data[9631] <= r_data[9630];
                
                r_data[9632] <= r_data[9631];
                
                r_data[9633] <= r_data[9632];
                
                r_data[9634] <= r_data[9633];
                
                r_data[9635] <= r_data[9634];
                
                r_data[9636] <= r_data[9635];
                
                r_data[9637] <= r_data[9636];
                
                r_data[9638] <= r_data[9637];
                
                r_data[9639] <= r_data[9638];
                
                r_data[9640] <= r_data[9639];
                
                r_data[9641] <= r_data[9640];
                
                r_data[9642] <= r_data[9641];
                
                r_data[9643] <= r_data[9642];
                
                r_data[9644] <= r_data[9643];
                
                r_data[9645] <= r_data[9644];
                
                r_data[9646] <= r_data[9645];
                
                r_data[9647] <= r_data[9646];
                
                r_data[9648] <= r_data[9647];
                
                r_data[9649] <= r_data[9648];
                
                r_data[9650] <= r_data[9649];
                
                r_data[9651] <= r_data[9650];
                
                r_data[9652] <= r_data[9651];
                
                r_data[9653] <= r_data[9652];
                
                r_data[9654] <= r_data[9653];
                
                r_data[9655] <= r_data[9654];
                
                r_data[9656] <= r_data[9655];
                
                r_data[9657] <= r_data[9656];
                
                r_data[9658] <= r_data[9657];
                
                r_data[9659] <= r_data[9658];
                
                r_data[9660] <= r_data[9659];
                
                r_data[9661] <= r_data[9660];
                
                r_data[9662] <= r_data[9661];
                
                r_data[9663] <= r_data[9662];
                
                r_data[9664] <= r_data[9663];
                
                r_data[9665] <= r_data[9664];
                
                r_data[9666] <= r_data[9665];
                
                r_data[9667] <= r_data[9666];
                
                r_data[9668] <= r_data[9667];
                
                r_data[9669] <= r_data[9668];
                
                r_data[9670] <= r_data[9669];
                
                r_data[9671] <= r_data[9670];
                
                r_data[9672] <= r_data[9671];
                
                r_data[9673] <= r_data[9672];
                
                r_data[9674] <= r_data[9673];
                
                r_data[9675] <= r_data[9674];
                
                r_data[9676] <= r_data[9675];
                
                r_data[9677] <= r_data[9676];
                
                r_data[9678] <= r_data[9677];
                
                r_data[9679] <= r_data[9678];
                
                r_data[9680] <= r_data[9679];
                
                r_data[9681] <= r_data[9680];
                
                r_data[9682] <= r_data[9681];
                
                r_data[9683] <= r_data[9682];
                
                r_data[9684] <= r_data[9683];
                
                r_data[9685] <= r_data[9684];
                
                r_data[9686] <= r_data[9685];
                
                r_data[9687] <= r_data[9686];
                
                r_data[9688] <= r_data[9687];
                
                r_data[9689] <= r_data[9688];
                
                r_data[9690] <= r_data[9689];
                
                r_data[9691] <= r_data[9690];
                
                r_data[9692] <= r_data[9691];
                
                r_data[9693] <= r_data[9692];
                
                r_data[9694] <= r_data[9693];
                
                r_data[9695] <= r_data[9694];
                
                r_data[9696] <= r_data[9695];
                
                r_data[9697] <= r_data[9696];
                
                r_data[9698] <= r_data[9697];
                
                r_data[9699] <= r_data[9698];
                
                r_data[9700] <= r_data[9699];
                
                r_data[9701] <= r_data[9700];
                
                r_data[9702] <= r_data[9701];
                
                r_data[9703] <= r_data[9702];
                
                r_data[9704] <= r_data[9703];
                
                r_data[9705] <= r_data[9704];
                
                r_data[9706] <= r_data[9705];
                
                r_data[9707] <= r_data[9706];
                
                r_data[9708] <= r_data[9707];
                
                r_data[9709] <= r_data[9708];
                
                r_data[9710] <= r_data[9709];
                
                r_data[9711] <= r_data[9710];
                
                r_data[9712] <= r_data[9711];
                
                r_data[9713] <= r_data[9712];
                
                r_data[9714] <= r_data[9713];
                
                r_data[9715] <= r_data[9714];
                
                r_data[9716] <= r_data[9715];
                
                r_data[9717] <= r_data[9716];
                
                r_data[9718] <= r_data[9717];
                
                r_data[9719] <= r_data[9718];
                
                r_data[9720] <= r_data[9719];
                
                r_data[9721] <= r_data[9720];
                
                r_data[9722] <= r_data[9721];
                
                r_data[9723] <= r_data[9722];
                
                r_data[9724] <= r_data[9723];
                
                r_data[9725] <= r_data[9724];
                
                r_data[9726] <= r_data[9725];
                
                r_data[9727] <= r_data[9726];
                
                r_data[9728] <= r_data[9727];
                
                r_data[9729] <= r_data[9728];
                
                r_data[9730] <= r_data[9729];
                
                r_data[9731] <= r_data[9730];
                
                r_data[9732] <= r_data[9731];
                
                r_data[9733] <= r_data[9732];
                
                r_data[9734] <= r_data[9733];
                
                r_data[9735] <= r_data[9734];
                
                r_data[9736] <= r_data[9735];
                
                r_data[9737] <= r_data[9736];
                
                r_data[9738] <= r_data[9737];
                
                r_data[9739] <= r_data[9738];
                
                r_data[9740] <= r_data[9739];
                
                r_data[9741] <= r_data[9740];
                
                r_data[9742] <= r_data[9741];
                
                r_data[9743] <= r_data[9742];
                
                r_data[9744] <= r_data[9743];
                
                r_data[9745] <= r_data[9744];
                
                r_data[9746] <= r_data[9745];
                
                r_data[9747] <= r_data[9746];
                
                r_data[9748] <= r_data[9747];
                
                r_data[9749] <= r_data[9748];
                
                r_data[9750] <= r_data[9749];
                
                r_data[9751] <= r_data[9750];
                
                r_data[9752] <= r_data[9751];
                
                r_data[9753] <= r_data[9752];
                
                r_data[9754] <= r_data[9753];
                
                r_data[9755] <= r_data[9754];
                
                r_data[9756] <= r_data[9755];
                
                r_data[9757] <= r_data[9756];
                
                r_data[9758] <= r_data[9757];
                
                r_data[9759] <= r_data[9758];
                
                r_data[9760] <= r_data[9759];
                
                r_data[9761] <= r_data[9760];
                
                r_data[9762] <= r_data[9761];
                
                r_data[9763] <= r_data[9762];
                
                r_data[9764] <= r_data[9763];
                
                r_data[9765] <= r_data[9764];
                
                r_data[9766] <= r_data[9765];
                
                r_data[9767] <= r_data[9766];
                
                r_data[9768] <= r_data[9767];
                
                r_data[9769] <= r_data[9768];
                
                r_data[9770] <= r_data[9769];
                
                r_data[9771] <= r_data[9770];
                
                r_data[9772] <= r_data[9771];
                
                r_data[9773] <= r_data[9772];
                
                r_data[9774] <= r_data[9773];
                
                r_data[9775] <= r_data[9774];
                
                r_data[9776] <= r_data[9775];
                
                r_data[9777] <= r_data[9776];
                
                r_data[9778] <= r_data[9777];
                
                r_data[9779] <= r_data[9778];
                
                r_data[9780] <= r_data[9779];
                
                r_data[9781] <= r_data[9780];
                
                r_data[9782] <= r_data[9781];
                
                r_data[9783] <= r_data[9782];
                
                r_data[9784] <= r_data[9783];
                
                r_data[9785] <= r_data[9784];
                
                r_data[9786] <= r_data[9785];
                
                r_data[9787] <= r_data[9786];
                
                r_data[9788] <= r_data[9787];
                
                r_data[9789] <= r_data[9788];
                
                r_data[9790] <= r_data[9789];
                
                r_data[9791] <= r_data[9790];
                
                r_data[9792] <= r_data[9791];
                
                r_data[9793] <= r_data[9792];
                
                r_data[9794] <= r_data[9793];
                
                r_data[9795] <= r_data[9794];
                
                r_data[9796] <= r_data[9795];
                
                r_data[9797] <= r_data[9796];
                
                r_data[9798] <= r_data[9797];
                
                r_data[9799] <= r_data[9798];
                
                r_data[9800] <= r_data[9799];
                
                r_data[9801] <= r_data[9800];
                
                r_data[9802] <= r_data[9801];
                
                r_data[9803] <= r_data[9802];
                
                r_data[9804] <= r_data[9803];
                
                r_data[9805] <= r_data[9804];
                
                r_data[9806] <= r_data[9805];
                
                r_data[9807] <= r_data[9806];
                
                r_data[9808] <= r_data[9807];
                
                r_data[9809] <= r_data[9808];
                
                r_data[9810] <= r_data[9809];
                
                r_data[9811] <= r_data[9810];
                
                r_data[9812] <= r_data[9811];
                
                r_data[9813] <= r_data[9812];
                
                r_data[9814] <= r_data[9813];
                
                r_data[9815] <= r_data[9814];
                
                r_data[9816] <= r_data[9815];
                
                r_data[9817] <= r_data[9816];
                
                r_data[9818] <= r_data[9817];
                
                r_data[9819] <= r_data[9818];
                
                r_data[9820] <= r_data[9819];
                
                r_data[9821] <= r_data[9820];
                
                r_data[9822] <= r_data[9821];
                
                r_data[9823] <= r_data[9822];
                
                r_data[9824] <= r_data[9823];
                
                r_data[9825] <= r_data[9824];
                
                r_data[9826] <= r_data[9825];
                
                r_data[9827] <= r_data[9826];
                
                r_data[9828] <= r_data[9827];
                
                r_data[9829] <= r_data[9828];
                
                r_data[9830] <= r_data[9829];
                
                r_data[9831] <= r_data[9830];
                
                r_data[9832] <= r_data[9831];
                
                r_data[9833] <= r_data[9832];
                
                r_data[9834] <= r_data[9833];
                
                r_data[9835] <= r_data[9834];
                
                r_data[9836] <= r_data[9835];
                
                r_data[9837] <= r_data[9836];
                
                r_data[9838] <= r_data[9837];
                
                r_data[9839] <= r_data[9838];
                
                r_data[9840] <= r_data[9839];
                
                r_data[9841] <= r_data[9840];
                
                r_data[9842] <= r_data[9841];
                
                r_data[9843] <= r_data[9842];
                
                r_data[9844] <= r_data[9843];
                
                r_data[9845] <= r_data[9844];
                
                r_data[9846] <= r_data[9845];
                
                r_data[9847] <= r_data[9846];
                
                r_data[9848] <= r_data[9847];
                
                r_data[9849] <= r_data[9848];
                
                r_data[9850] <= r_data[9849];
                
                r_data[9851] <= r_data[9850];
                
                r_data[9852] <= r_data[9851];
                
                r_data[9853] <= r_data[9852];
                
                r_data[9854] <= r_data[9853];
                
                r_data[9855] <= r_data[9854];
                
                r_data[9856] <= r_data[9855];
                
                r_data[9857] <= r_data[9856];
                
                r_data[9858] <= r_data[9857];
                
                r_data[9859] <= r_data[9858];
                
                r_data[9860] <= r_data[9859];
                
                r_data[9861] <= r_data[9860];
                
                r_data[9862] <= r_data[9861];
                
                r_data[9863] <= r_data[9862];
                
                r_data[9864] <= r_data[9863];
                
                r_data[9865] <= r_data[9864];
                
                r_data[9866] <= r_data[9865];
                
                r_data[9867] <= r_data[9866];
                
                r_data[9868] <= r_data[9867];
                
                r_data[9869] <= r_data[9868];
                
                r_data[9870] <= r_data[9869];
                
                r_data[9871] <= r_data[9870];
                
                r_data[9872] <= r_data[9871];
                
                r_data[9873] <= r_data[9872];
                
                r_data[9874] <= r_data[9873];
                
                r_data[9875] <= r_data[9874];
                
                r_data[9876] <= r_data[9875];
                
                r_data[9877] <= r_data[9876];
                
                r_data[9878] <= r_data[9877];
                
                r_data[9879] <= r_data[9878];
                
                r_data[9880] <= r_data[9879];
                
                r_data[9881] <= r_data[9880];
                
                r_data[9882] <= r_data[9881];
                
                r_data[9883] <= r_data[9882];
                
                r_data[9884] <= r_data[9883];
                
                r_data[9885] <= r_data[9884];
                
                r_data[9886] <= r_data[9885];
                
                r_data[9887] <= r_data[9886];
                
                r_data[9888] <= r_data[9887];
                
                r_data[9889] <= r_data[9888];
                
                r_data[9890] <= r_data[9889];
                
                r_data[9891] <= r_data[9890];
                
                r_data[9892] <= r_data[9891];
                
                r_data[9893] <= r_data[9892];
                
                r_data[9894] <= r_data[9893];
                
                r_data[9895] <= r_data[9894];
                
                r_data[9896] <= r_data[9895];
                
                r_data[9897] <= r_data[9896];
                
                r_data[9898] <= r_data[9897];
                
                r_data[9899] <= r_data[9898];
                
                r_data[9900] <= r_data[9899];
                
                r_data[9901] <= r_data[9900];
                
                r_data[9902] <= r_data[9901];
                
                r_data[9903] <= r_data[9902];
                
                r_data[9904] <= r_data[9903];
                
                r_data[9905] <= r_data[9904];
                
                r_data[9906] <= r_data[9905];
                
                r_data[9907] <= r_data[9906];
                
                r_data[9908] <= r_data[9907];
                
                r_data[9909] <= r_data[9908];
                
                r_data[9910] <= r_data[9909];
                
                r_data[9911] <= r_data[9910];
                
                r_data[9912] <= r_data[9911];
                
                r_data[9913] <= r_data[9912];
                
                r_data[9914] <= r_data[9913];
                
                r_data[9915] <= r_data[9914];
                
                r_data[9916] <= r_data[9915];
                
                r_data[9917] <= r_data[9916];
                
                r_data[9918] <= r_data[9917];
                
                r_data[9919] <= r_data[9918];
                
                r_data[9920] <= r_data[9919];
                
                r_data[9921] <= r_data[9920];
                
                r_data[9922] <= r_data[9921];
                
                r_data[9923] <= r_data[9922];
                
                r_data[9924] <= r_data[9923];
                
                r_data[9925] <= r_data[9924];
                
                r_data[9926] <= r_data[9925];
                
                r_data[9927] <= r_data[9926];
                
                r_data[9928] <= r_data[9927];
                
                r_data[9929] <= r_data[9928];
                
                r_data[9930] <= r_data[9929];
                
                r_data[9931] <= r_data[9930];
                
                r_data[9932] <= r_data[9931];
                
                r_data[9933] <= r_data[9932];
                
                r_data[9934] <= r_data[9933];
                
                r_data[9935] <= r_data[9934];
                
                r_data[9936] <= r_data[9935];
                
                r_data[9937] <= r_data[9936];
                
                r_data[9938] <= r_data[9937];
                
                r_data[9939] <= r_data[9938];
                
                r_data[9940] <= r_data[9939];
                
                r_data[9941] <= r_data[9940];
                
                r_data[9942] <= r_data[9941];
                
                r_data[9943] <= r_data[9942];
                
                r_data[9944] <= r_data[9943];
                
                r_data[9945] <= r_data[9944];
                
                r_data[9946] <= r_data[9945];
                
                r_data[9947] <= r_data[9946];
                
                r_data[9948] <= r_data[9947];
                
                r_data[9949] <= r_data[9948];
                
                r_data[9950] <= r_data[9949];
                
                r_data[9951] <= r_data[9950];
                
                r_data[9952] <= r_data[9951];
                
                r_data[9953] <= r_data[9952];
                
                r_data[9954] <= r_data[9953];
                
                r_data[9955] <= r_data[9954];
                
                r_data[9956] <= r_data[9955];
                
                r_data[9957] <= r_data[9956];
                
                r_data[9958] <= r_data[9957];
                
                r_data[9959] <= r_data[9958];
                
                r_data[9960] <= r_data[9959];
                
                r_data[9961] <= r_data[9960];
                
                r_data[9962] <= r_data[9961];
                
                r_data[9963] <= r_data[9962];
                
                r_data[9964] <= r_data[9963];
                
                r_data[9965] <= r_data[9964];
                
                r_data[9966] <= r_data[9965];
                
                r_data[9967] <= r_data[9966];
                
                r_data[9968] <= r_data[9967];
                
                r_data[9969] <= r_data[9968];
                
                r_data[9970] <= r_data[9969];
                
                r_data[9971] <= r_data[9970];
                
                r_data[9972] <= r_data[9971];
                
                r_data[9973] <= r_data[9972];
                
                r_data[9974] <= r_data[9973];
                
                r_data[9975] <= r_data[9974];
                
                r_data[9976] <= r_data[9975];
                
                r_data[9977] <= r_data[9976];
                
                r_data[9978] <= r_data[9977];
                
                r_data[9979] <= r_data[9978];
                
                r_data[9980] <= r_data[9979];
                
                r_data[9981] <= r_data[9980];
                
                r_data[9982] <= r_data[9981];
                
                r_data[9983] <= r_data[9982];
                
                r_data[9984] <= r_data[9983];
                
                r_data[9985] <= r_data[9984];
                
                r_data[9986] <= r_data[9985];
                
                r_data[9987] <= r_data[9986];
                
                r_data[9988] <= r_data[9987];
                
                r_data[9989] <= r_data[9988];
                
                r_data[9990] <= r_data[9989];
                
                r_data[9991] <= r_data[9990];
                
                r_data[9992] <= r_data[9991];
                
                r_data[9993] <= r_data[9992];
                
                r_data[9994] <= r_data[9993];
                
                r_data[9995] <= r_data[9994];
                
                r_data[9996] <= r_data[9995];
                
                r_data[9997] <= r_data[9996];
                
                r_data[9998] <= r_data[9997];
                
                r_data[9999] <= r_data[9998];
                
                r_data[10000] <= r_data[9999];
                
                r_data[10001] <= r_data[10000];
                
                r_data[10002] <= r_data[10001];
                
                r_data[10003] <= r_data[10002];
                
                r_data[10004] <= r_data[10003];
                
                r_data[10005] <= r_data[10004];
                
                r_data[10006] <= r_data[10005];
                
                r_data[10007] <= r_data[10006];
                
                r_data[10008] <= r_data[10007];
                
                r_data[10009] <= r_data[10008];
                
                r_data[10010] <= r_data[10009];
                
                r_data[10011] <= r_data[10010];
                
                r_data[10012] <= r_data[10011];
                
                r_data[10013] <= r_data[10012];
                
                r_data[10014] <= r_data[10013];
                
                r_data[10015] <= r_data[10014];
                
                r_data[10016] <= r_data[10015];
                
                r_data[10017] <= r_data[10016];
                
                r_data[10018] <= r_data[10017];
                
                r_data[10019] <= r_data[10018];
                
                r_data[10020] <= r_data[10019];
                
                r_data[10021] <= r_data[10020];
                
                r_data[10022] <= r_data[10021];
                
                r_data[10023] <= r_data[10022];
                
                r_data[10024] <= r_data[10023];
                
                r_data[10025] <= r_data[10024];
                
                r_data[10026] <= r_data[10025];
                
                r_data[10027] <= r_data[10026];
                
                r_data[10028] <= r_data[10027];
                
                r_data[10029] <= r_data[10028];
                
                r_data[10030] <= r_data[10029];
                
                r_data[10031] <= r_data[10030];
                
                r_data[10032] <= r_data[10031];
                
                r_data[10033] <= r_data[10032];
                
                r_data[10034] <= r_data[10033];
                
                r_data[10035] <= r_data[10034];
                
                r_data[10036] <= r_data[10035];
                
                r_data[10037] <= r_data[10036];
                
                r_data[10038] <= r_data[10037];
                
                r_data[10039] <= r_data[10038];
                
                r_data[10040] <= r_data[10039];
                
                r_data[10041] <= r_data[10040];
                
                r_data[10042] <= r_data[10041];
                
                r_data[10043] <= r_data[10042];
                
                r_data[10044] <= r_data[10043];
                
                r_data[10045] <= r_data[10044];
                
                r_data[10046] <= r_data[10045];
                
                r_data[10047] <= r_data[10046];
                
                r_data[10048] <= r_data[10047];
                
                r_data[10049] <= r_data[10048];
                
                r_data[10050] <= r_data[10049];
                
                r_data[10051] <= r_data[10050];
                
                r_data[10052] <= r_data[10051];
                
                r_data[10053] <= r_data[10052];
                
                r_data[10054] <= r_data[10053];
                
                r_data[10055] <= r_data[10054];
                
                r_data[10056] <= r_data[10055];
                
                r_data[10057] <= r_data[10056];
                
                r_data[10058] <= r_data[10057];
                
                r_data[10059] <= r_data[10058];
                
                r_data[10060] <= r_data[10059];
                
                r_data[10061] <= r_data[10060];
                
                r_data[10062] <= r_data[10061];
                
                r_data[10063] <= r_data[10062];
                
                r_data[10064] <= r_data[10063];
                
                r_data[10065] <= r_data[10064];
                
                r_data[10066] <= r_data[10065];
                
                r_data[10067] <= r_data[10066];
                
                r_data[10068] <= r_data[10067];
                
                r_data[10069] <= r_data[10068];
                
                r_data[10070] <= r_data[10069];
                
                r_data[10071] <= r_data[10070];
                
                r_data[10072] <= r_data[10071];
                
                r_data[10073] <= r_data[10072];
                
                r_data[10074] <= r_data[10073];
                
                r_data[10075] <= r_data[10074];
                
                r_data[10076] <= r_data[10075];
                
                r_data[10077] <= r_data[10076];
                
                r_data[10078] <= r_data[10077];
                
                r_data[10079] <= r_data[10078];
                
                r_data[10080] <= r_data[10079];
                
                r_data[10081] <= r_data[10080];
                
                r_data[10082] <= r_data[10081];
                
                r_data[10083] <= r_data[10082];
                
                r_data[10084] <= r_data[10083];
                
                r_data[10085] <= r_data[10084];
                
                r_data[10086] <= r_data[10085];
                
                r_data[10087] <= r_data[10086];
                
                r_data[10088] <= r_data[10087];
                
                r_data[10089] <= r_data[10088];
                
                r_data[10090] <= r_data[10089];
                
                r_data[10091] <= r_data[10090];
                
                r_data[10092] <= r_data[10091];
                
                r_data[10093] <= r_data[10092];
                
                r_data[10094] <= r_data[10093];
                
                r_data[10095] <= r_data[10094];
                
                r_data[10096] <= r_data[10095];
                
                r_data[10097] <= r_data[10096];
                
                r_data[10098] <= r_data[10097];
                
                r_data[10099] <= r_data[10098];
                
                r_data[10100] <= r_data[10099];
                
                r_data[10101] <= r_data[10100];
                
                r_data[10102] <= r_data[10101];
                
                r_data[10103] <= r_data[10102];
                
                r_data[10104] <= r_data[10103];
                
                r_data[10105] <= r_data[10104];
                
                r_data[10106] <= r_data[10105];
                
                r_data[10107] <= r_data[10106];
                
                r_data[10108] <= r_data[10107];
                
                r_data[10109] <= r_data[10108];
                
                r_data[10110] <= r_data[10109];
                
                r_data[10111] <= r_data[10110];
                
                r_data[10112] <= r_data[10111];
                
                r_data[10113] <= r_data[10112];
                
                r_data[10114] <= r_data[10113];
                
                r_data[10115] <= r_data[10114];
                
                r_data[10116] <= r_data[10115];
                
                r_data[10117] <= r_data[10116];
                
                r_data[10118] <= r_data[10117];
                
                r_data[10119] <= r_data[10118];
                
                r_data[10120] <= r_data[10119];
                
                r_data[10121] <= r_data[10120];
                
                r_data[10122] <= r_data[10121];
                
                r_data[10123] <= r_data[10122];
                
                r_data[10124] <= r_data[10123];
                
                r_data[10125] <= r_data[10124];
                
                r_data[10126] <= r_data[10125];
                
                r_data[10127] <= r_data[10126];
                
                r_data[10128] <= r_data[10127];
                
                r_data[10129] <= r_data[10128];
                
                r_data[10130] <= r_data[10129];
                
                r_data[10131] <= r_data[10130];
                
                r_data[10132] <= r_data[10131];
                
                r_data[10133] <= r_data[10132];
                
                r_data[10134] <= r_data[10133];
                
                r_data[10135] <= r_data[10134];
                
                r_data[10136] <= r_data[10135];
                
                r_data[10137] <= r_data[10136];
                
                r_data[10138] <= r_data[10137];
                
                r_data[10139] <= r_data[10138];
                
                r_data[10140] <= r_data[10139];
                
                r_data[10141] <= r_data[10140];
                
                r_data[10142] <= r_data[10141];
                
                r_data[10143] <= r_data[10142];
                
                r_data[10144] <= r_data[10143];
                
                r_data[10145] <= r_data[10144];
                
                r_data[10146] <= r_data[10145];
                
                r_data[10147] <= r_data[10146];
                
                r_data[10148] <= r_data[10147];
                
                r_data[10149] <= r_data[10148];
                
                r_data[10150] <= r_data[10149];
                
                r_data[10151] <= r_data[10150];
                
                r_data[10152] <= r_data[10151];
                
                r_data[10153] <= r_data[10152];
                
                r_data[10154] <= r_data[10153];
                
                r_data[10155] <= r_data[10154];
                
                r_data[10156] <= r_data[10155];
                
                r_data[10157] <= r_data[10156];
                
                r_data[10158] <= r_data[10157];
                
                r_data[10159] <= r_data[10158];
                
                r_data[10160] <= r_data[10159];
                
                r_data[10161] <= r_data[10160];
                
                r_data[10162] <= r_data[10161];
                
                r_data[10163] <= r_data[10162];
                
                r_data[10164] <= r_data[10163];
                
                r_data[10165] <= r_data[10164];
                
                r_data[10166] <= r_data[10165];
                
                r_data[10167] <= r_data[10166];
                
                r_data[10168] <= r_data[10167];
                
                r_data[10169] <= r_data[10168];
                
                r_data[10170] <= r_data[10169];
                
                r_data[10171] <= r_data[10170];
                
                r_data[10172] <= r_data[10171];
                
                r_data[10173] <= r_data[10172];
                
                r_data[10174] <= r_data[10173];
                
                r_data[10175] <= r_data[10174];
                
                r_data[10176] <= r_data[10175];
                
                r_data[10177] <= r_data[10176];
                
                r_data[10178] <= r_data[10177];
                
                r_data[10179] <= r_data[10178];
                
                r_data[10180] <= r_data[10179];
                
                r_data[10181] <= r_data[10180];
                
                r_data[10182] <= r_data[10181];
                
                r_data[10183] <= r_data[10182];
                
                r_data[10184] <= r_data[10183];
                
                r_data[10185] <= r_data[10184];
                
                r_data[10186] <= r_data[10185];
                
                r_data[10187] <= r_data[10186];
                
                r_data[10188] <= r_data[10187];
                
                r_data[10189] <= r_data[10188];
                
                r_data[10190] <= r_data[10189];
                
                r_data[10191] <= r_data[10190];
                
                r_data[10192] <= r_data[10191];
                
                r_data[10193] <= r_data[10192];
                
                r_data[10194] <= r_data[10193];
                
                r_data[10195] <= r_data[10194];
                
                r_data[10196] <= r_data[10195];
                
                r_data[10197] <= r_data[10196];
                
                r_data[10198] <= r_data[10197];
                
                r_data[10199] <= r_data[10198];
                
                r_data[10200] <= r_data[10199];
                
                r_data[10201] <= r_data[10200];
                
                r_data[10202] <= r_data[10201];
                
                r_data[10203] <= r_data[10202];
                
                r_data[10204] <= r_data[10203];
                
                r_data[10205] <= r_data[10204];
                
                r_data[10206] <= r_data[10205];
                
                r_data[10207] <= r_data[10206];
                
                r_data[10208] <= r_data[10207];
                
                r_data[10209] <= r_data[10208];
                
                r_data[10210] <= r_data[10209];
                
                r_data[10211] <= r_data[10210];
                
                r_data[10212] <= r_data[10211];
                
                r_data[10213] <= r_data[10212];
                
                r_data[10214] <= r_data[10213];
                
                r_data[10215] <= r_data[10214];
                
                r_data[10216] <= r_data[10215];
                
                r_data[10217] <= r_data[10216];
                
                r_data[10218] <= r_data[10217];
                
                r_data[10219] <= r_data[10218];
                
                r_data[10220] <= r_data[10219];
                
                r_data[10221] <= r_data[10220];
                
                r_data[10222] <= r_data[10221];
                
                r_data[10223] <= r_data[10222];
                
                r_data[10224] <= r_data[10223];
                
                r_data[10225] <= r_data[10224];
                
                r_data[10226] <= r_data[10225];
                
                r_data[10227] <= r_data[10226];
                
                r_data[10228] <= r_data[10227];
                
                r_data[10229] <= r_data[10228];
                
                r_data[10230] <= r_data[10229];
                
                r_data[10231] <= r_data[10230];
                
                r_data[10232] <= r_data[10231];
                
                r_data[10233] <= r_data[10232];
                
                r_data[10234] <= r_data[10233];
                
                r_data[10235] <= r_data[10234];
                
                r_data[10236] <= r_data[10235];
                
                r_data[10237] <= r_data[10236];
                
                r_data[10238] <= r_data[10237];
                
                r_data[10239] <= r_data[10238];
                
                r_data[10240] <= r_data[10239];
                
                r_data[10241] <= r_data[10240];
                
                r_data[10242] <= r_data[10241];
                
                r_data[10243] <= r_data[10242];
                
                r_data[10244] <= r_data[10243];
                
                r_data[10245] <= r_data[10244];
                
                r_data[10246] <= r_data[10245];
                
                r_data[10247] <= r_data[10246];
                
                r_data[10248] <= r_data[10247];
                
                r_data[10249] <= r_data[10248];
                
                r_data[10250] <= r_data[10249];
                
                r_data[10251] <= r_data[10250];
                
                r_data[10252] <= r_data[10251];
                
                r_data[10253] <= r_data[10252];
                
                r_data[10254] <= r_data[10253];
                
                r_data[10255] <= r_data[10254];
                
                r_data[10256] <= r_data[10255];
                
                r_data[10257] <= r_data[10256];
                
                r_data[10258] <= r_data[10257];
                
                r_data[10259] <= r_data[10258];
                
                r_data[10260] <= r_data[10259];
                
                r_data[10261] <= r_data[10260];
                
                r_data[10262] <= r_data[10261];
                
                r_data[10263] <= r_data[10262];
                
                r_data[10264] <= r_data[10263];
                
                r_data[10265] <= r_data[10264];
                
                r_data[10266] <= r_data[10265];
                
                r_data[10267] <= r_data[10266];
                
                r_data[10268] <= r_data[10267];
                
                r_data[10269] <= r_data[10268];
                
                r_data[10270] <= r_data[10269];
                
                r_data[10271] <= r_data[10270];
                
                r_data[10272] <= r_data[10271];
                
                r_data[10273] <= r_data[10272];
                
                r_data[10274] <= r_data[10273];
                
                r_data[10275] <= r_data[10274];
                
                r_data[10276] <= r_data[10275];
                
                r_data[10277] <= r_data[10276];
                
                r_data[10278] <= r_data[10277];
                
                r_data[10279] <= r_data[10278];
                
                r_data[10280] <= r_data[10279];
                
                r_data[10281] <= r_data[10280];
                
                r_data[10282] <= r_data[10281];
                
                r_data[10283] <= r_data[10282];
                
                r_data[10284] <= r_data[10283];
                
                r_data[10285] <= r_data[10284];
                
                r_data[10286] <= r_data[10285];
                
                r_data[10287] <= r_data[10286];
                
                r_data[10288] <= r_data[10287];
                
                r_data[10289] <= r_data[10288];
                
                r_data[10290] <= r_data[10289];
                
                r_data[10291] <= r_data[10290];
                
                r_data[10292] <= r_data[10291];
                
                r_data[10293] <= r_data[10292];
                
                r_data[10294] <= r_data[10293];
                
                r_data[10295] <= r_data[10294];
                
                r_data[10296] <= r_data[10295];
                
                r_data[10297] <= r_data[10296];
                
                r_data[10298] <= r_data[10297];
                
                r_data[10299] <= r_data[10298];
                
                r_data[10300] <= r_data[10299];
                
                r_data[10301] <= r_data[10300];
                
                r_data[10302] <= r_data[10301];
                
                r_data[10303] <= r_data[10302];
                
                r_data[10304] <= r_data[10303];
                
                r_data[10305] <= r_data[10304];
                
                r_data[10306] <= r_data[10305];
                
                r_data[10307] <= r_data[10306];
                
                r_data[10308] <= r_data[10307];
                
                r_data[10309] <= r_data[10308];
                
                r_data[10310] <= r_data[10309];
                
                r_data[10311] <= r_data[10310];
                
                r_data[10312] <= r_data[10311];
                
                r_data[10313] <= r_data[10312];
                
                r_data[10314] <= r_data[10313];
                
                r_data[10315] <= r_data[10314];
                
                r_data[10316] <= r_data[10315];
                
                r_data[10317] <= r_data[10316];
                
                r_data[10318] <= r_data[10317];
                
                r_data[10319] <= r_data[10318];
                
                r_data[10320] <= r_data[10319];
                
                r_data[10321] <= r_data[10320];
                
                r_data[10322] <= r_data[10321];
                
                r_data[10323] <= r_data[10322];
                
                r_data[10324] <= r_data[10323];
                
                r_data[10325] <= r_data[10324];
                
                r_data[10326] <= r_data[10325];
                
                r_data[10327] <= r_data[10326];
                
                r_data[10328] <= r_data[10327];
                
                r_data[10329] <= r_data[10328];
                
                r_data[10330] <= r_data[10329];
                
                r_data[10331] <= r_data[10330];
                
                r_data[10332] <= r_data[10331];
                
                r_data[10333] <= r_data[10332];
                
                r_data[10334] <= r_data[10333];
                
                r_data[10335] <= r_data[10334];
                
                r_data[10336] <= r_data[10335];
                
                r_data[10337] <= r_data[10336];
                
                r_data[10338] <= r_data[10337];
                
                r_data[10339] <= r_data[10338];
                
                r_data[10340] <= r_data[10339];
                
                r_data[10341] <= r_data[10340];
                
                r_data[10342] <= r_data[10341];
                
                r_data[10343] <= r_data[10342];
                
                r_data[10344] <= r_data[10343];
                
                r_data[10345] <= r_data[10344];
                
                r_data[10346] <= r_data[10345];
                
                r_data[10347] <= r_data[10346];
                
                r_data[10348] <= r_data[10347];
                
                r_data[10349] <= r_data[10348];
                
                r_data[10350] <= r_data[10349];
                
                r_data[10351] <= r_data[10350];
                
                r_data[10352] <= r_data[10351];
                
                r_data[10353] <= r_data[10352];
                
                r_data[10354] <= r_data[10353];
                
                r_data[10355] <= r_data[10354];
                
                r_data[10356] <= r_data[10355];
                
                r_data[10357] <= r_data[10356];
                
                r_data[10358] <= r_data[10357];
                
                r_data[10359] <= r_data[10358];
                
                r_data[10360] <= r_data[10359];
                
                r_data[10361] <= r_data[10360];
                
                r_data[10362] <= r_data[10361];
                
                r_data[10363] <= r_data[10362];
                
                r_data[10364] <= r_data[10363];
                
                r_data[10365] <= r_data[10364];
                
                r_data[10366] <= r_data[10365];
                
                r_data[10367] <= r_data[10366];
                
                r_data[10368] <= r_data[10367];
                
                r_data[10369] <= r_data[10368];
                
                r_data[10370] <= r_data[10369];
                
                r_data[10371] <= r_data[10370];
                
                r_data[10372] <= r_data[10371];
                
                r_data[10373] <= r_data[10372];
                
                r_data[10374] <= r_data[10373];
                
                r_data[10375] <= r_data[10374];
                
                r_data[10376] <= r_data[10375];
                
                r_data[10377] <= r_data[10376];
                
                r_data[10378] <= r_data[10377];
                
                r_data[10379] <= r_data[10378];
                
                r_data[10380] <= r_data[10379];
                
                r_data[10381] <= r_data[10380];
                
                r_data[10382] <= r_data[10381];
                
                r_data[10383] <= r_data[10382];
                
                r_data[10384] <= r_data[10383];
                
                r_data[10385] <= r_data[10384];
                
                r_data[10386] <= r_data[10385];
                
                r_data[10387] <= r_data[10386];
                
                r_data[10388] <= r_data[10387];
                
                r_data[10389] <= r_data[10388];
                
                r_data[10390] <= r_data[10389];
                
                r_data[10391] <= r_data[10390];
                
                r_data[10392] <= r_data[10391];
                
                r_data[10393] <= r_data[10392];
                
                r_data[10394] <= r_data[10393];
                
                r_data[10395] <= r_data[10394];
                
                r_data[10396] <= r_data[10395];
                
                r_data[10397] <= r_data[10396];
                
                r_data[10398] <= r_data[10397];
                
                r_data[10399] <= r_data[10398];
                
                r_data[10400] <= r_data[10399];
                
                r_data[10401] <= r_data[10400];
                
                r_data[10402] <= r_data[10401];
                
                r_data[10403] <= r_data[10402];
                
                r_data[10404] <= r_data[10403];
                
                r_data[10405] <= r_data[10404];
                
                r_data[10406] <= r_data[10405];
                
                r_data[10407] <= r_data[10406];
                
                r_data[10408] <= r_data[10407];
                
                r_data[10409] <= r_data[10408];
                
                r_data[10410] <= r_data[10409];
                
                r_data[10411] <= r_data[10410];
                
                r_data[10412] <= r_data[10411];
                
                r_data[10413] <= r_data[10412];
                
                r_data[10414] <= r_data[10413];
                
                r_data[10415] <= r_data[10414];
                
                r_data[10416] <= r_data[10415];
                
                r_data[10417] <= r_data[10416];
                
                r_data[10418] <= r_data[10417];
                
                r_data[10419] <= r_data[10418];
                
                r_data[10420] <= r_data[10419];
                
                r_data[10421] <= r_data[10420];
                
                r_data[10422] <= r_data[10421];
                
                r_data[10423] <= r_data[10422];
                
                r_data[10424] <= r_data[10423];
                
                r_data[10425] <= r_data[10424];
                
                r_data[10426] <= r_data[10425];
                
                r_data[10427] <= r_data[10426];
                
                r_data[10428] <= r_data[10427];
                
                r_data[10429] <= r_data[10428];
                
                r_data[10430] <= r_data[10429];
                
                r_data[10431] <= r_data[10430];
                
                r_data[10432] <= r_data[10431];
                
                r_data[10433] <= r_data[10432];
                
                r_data[10434] <= r_data[10433];
                
                r_data[10435] <= r_data[10434];
                
                r_data[10436] <= r_data[10435];
                
                r_data[10437] <= r_data[10436];
                
                r_data[10438] <= r_data[10437];
                
                r_data[10439] <= r_data[10438];
                
                r_data[10440] <= r_data[10439];
                
                r_data[10441] <= r_data[10440];
                
                r_data[10442] <= r_data[10441];
                
                r_data[10443] <= r_data[10442];
                
                r_data[10444] <= r_data[10443];
                
                r_data[10445] <= r_data[10444];
                
                r_data[10446] <= r_data[10445];
                
                r_data[10447] <= r_data[10446];
                
                r_data[10448] <= r_data[10447];
                
                r_data[10449] <= r_data[10448];
                
                r_data[10450] <= r_data[10449];
                
                r_data[10451] <= r_data[10450];
                
                r_data[10452] <= r_data[10451];
                
                r_data[10453] <= r_data[10452];
                
                r_data[10454] <= r_data[10453];
                
                r_data[10455] <= r_data[10454];
                
                r_data[10456] <= r_data[10455];
                
                r_data[10457] <= r_data[10456];
                
                r_data[10458] <= r_data[10457];
                
                r_data[10459] <= r_data[10458];
                
                r_data[10460] <= r_data[10459];
                
                r_data[10461] <= r_data[10460];
                
                r_data[10462] <= r_data[10461];
                
                r_data[10463] <= r_data[10462];
                
                r_data[10464] <= r_data[10463];
                
                r_data[10465] <= r_data[10464];
                
                r_data[10466] <= r_data[10465];
                
                r_data[10467] <= r_data[10466];
                
                r_data[10468] <= r_data[10467];
                
                r_data[10469] <= r_data[10468];
                
                r_data[10470] <= r_data[10469];
                
                r_data[10471] <= r_data[10470];
                
                r_data[10472] <= r_data[10471];
                
                r_data[10473] <= r_data[10472];
                
                r_data[10474] <= r_data[10473];
                
                r_data[10475] <= r_data[10474];
                
                r_data[10476] <= r_data[10475];
                
                r_data[10477] <= r_data[10476];
                
                r_data[10478] <= r_data[10477];
                
                r_data[10479] <= r_data[10478];
                
                r_data[10480] <= r_data[10479];
                
                r_data[10481] <= r_data[10480];
                
                r_data[10482] <= r_data[10481];
                
                r_data[10483] <= r_data[10482];
                
                r_data[10484] <= r_data[10483];
                
                r_data[10485] <= r_data[10484];
                
                r_data[10486] <= r_data[10485];
                
                r_data[10487] <= r_data[10486];
                
                r_data[10488] <= r_data[10487];
                
                r_data[10489] <= r_data[10488];
                
                r_data[10490] <= r_data[10489];
                
                r_data[10491] <= r_data[10490];
                
                r_data[10492] <= r_data[10491];
                
                r_data[10493] <= r_data[10492];
                
                r_data[10494] <= r_data[10493];
                
                r_data[10495] <= r_data[10494];
                
                r_data[10496] <= r_data[10495];
                
                r_data[10497] <= r_data[10496];
                
                r_data[10498] <= r_data[10497];
                
                r_data[10499] <= r_data[10498];
                
                r_data[10500] <= r_data[10499];
                
                r_data[10501] <= r_data[10500];
                
                r_data[10502] <= r_data[10501];
                
                r_data[10503] <= r_data[10502];
                
                r_data[10504] <= r_data[10503];
                
                r_data[10505] <= r_data[10504];
                
                r_data[10506] <= r_data[10505];
                
                r_data[10507] <= r_data[10506];
                
                r_data[10508] <= r_data[10507];
                
                r_data[10509] <= r_data[10508];
                
                r_data[10510] <= r_data[10509];
                
                r_data[10511] <= r_data[10510];
                
                r_data[10512] <= r_data[10511];
                
                r_data[10513] <= r_data[10512];
                
                r_data[10514] <= r_data[10513];
                
                r_data[10515] <= r_data[10514];
                
                r_data[10516] <= r_data[10515];
                
                r_data[10517] <= r_data[10516];
                
                r_data[10518] <= r_data[10517];
                
                r_data[10519] <= r_data[10518];
                
                r_data[10520] <= r_data[10519];
                
                r_data[10521] <= r_data[10520];
                
                r_data[10522] <= r_data[10521];
                
                r_data[10523] <= r_data[10522];
                
                r_data[10524] <= r_data[10523];
                
                r_data[10525] <= r_data[10524];
                
                r_data[10526] <= r_data[10525];
                
                r_data[10527] <= r_data[10526];
                
                r_data[10528] <= r_data[10527];
                
                r_data[10529] <= r_data[10528];
                
                r_data[10530] <= r_data[10529];
                
                r_data[10531] <= r_data[10530];
                
                r_data[10532] <= r_data[10531];
                
                r_data[10533] <= r_data[10532];
                
                r_data[10534] <= r_data[10533];
                
                r_data[10535] <= r_data[10534];
                
                r_data[10536] <= r_data[10535];
                
                r_data[10537] <= r_data[10536];
                
                r_data[10538] <= r_data[10537];
                
                r_data[10539] <= r_data[10538];
                
                r_data[10540] <= r_data[10539];
                
                r_data[10541] <= r_data[10540];
                
                r_data[10542] <= r_data[10541];
                
                r_data[10543] <= r_data[10542];
                
                r_data[10544] <= r_data[10543];
                
                r_data[10545] <= r_data[10544];
                
                r_data[10546] <= r_data[10545];
                
                r_data[10547] <= r_data[10546];
                
                r_data[10548] <= r_data[10547];
                
                r_data[10549] <= r_data[10548];
                
                r_data[10550] <= r_data[10549];
                
                r_data[10551] <= r_data[10550];
                
                r_data[10552] <= r_data[10551];
                
                r_data[10553] <= r_data[10552];
                
                r_data[10554] <= r_data[10553];
                
                r_data[10555] <= r_data[10554];
                
                r_data[10556] <= r_data[10555];
                
                r_data[10557] <= r_data[10556];
                
                r_data[10558] <= r_data[10557];
                
                r_data[10559] <= r_data[10558];
                
                r_data[10560] <= r_data[10559];
                
                r_data[10561] <= r_data[10560];
                
                r_data[10562] <= r_data[10561];
                
                r_data[10563] <= r_data[10562];
                
                r_data[10564] <= r_data[10563];
                
                r_data[10565] <= r_data[10564];
                
                r_data[10566] <= r_data[10565];
                
                r_data[10567] <= r_data[10566];
                
                r_data[10568] <= r_data[10567];
                
                r_data[10569] <= r_data[10568];
                
                r_data[10570] <= r_data[10569];
                
                r_data[10571] <= r_data[10570];
                
                r_data[10572] <= r_data[10571];
                
                r_data[10573] <= r_data[10572];
                
                r_data[10574] <= r_data[10573];
                
                r_data[10575] <= r_data[10574];
                
                r_data[10576] <= r_data[10575];
                
                r_data[10577] <= r_data[10576];
                
                r_data[10578] <= r_data[10577];
                
                r_data[10579] <= r_data[10578];
                
                r_data[10580] <= r_data[10579];
                
                r_data[10581] <= r_data[10580];
                
                r_data[10582] <= r_data[10581];
                
                r_data[10583] <= r_data[10582];
                
                r_data[10584] <= r_data[10583];
                
                r_data[10585] <= r_data[10584];
                
                r_data[10586] <= r_data[10585];
                
                r_data[10587] <= r_data[10586];
                
                r_data[10588] <= r_data[10587];
                
                r_data[10589] <= r_data[10588];
                
                r_data[10590] <= r_data[10589];
                
                r_data[10591] <= r_data[10590];
                
                r_data[10592] <= r_data[10591];
                
                r_data[10593] <= r_data[10592];
                
                r_data[10594] <= r_data[10593];
                
                r_data[10595] <= r_data[10594];
                
                r_data[10596] <= r_data[10595];
                
                r_data[10597] <= r_data[10596];
                
                r_data[10598] <= r_data[10597];
                
                r_data[10599] <= r_data[10598];
                
                r_data[10600] <= r_data[10599];
                
                r_data[10601] <= r_data[10600];
                
                r_data[10602] <= r_data[10601];
                
                r_data[10603] <= r_data[10602];
                
                r_data[10604] <= r_data[10603];
                
                r_data[10605] <= r_data[10604];
                
                r_data[10606] <= r_data[10605];
                
                r_data[10607] <= r_data[10606];
                
                r_data[10608] <= r_data[10607];
                
                r_data[10609] <= r_data[10608];
                
                r_data[10610] <= r_data[10609];
                
                r_data[10611] <= r_data[10610];
                
                r_data[10612] <= r_data[10611];
                
                r_data[10613] <= r_data[10612];
                
                r_data[10614] <= r_data[10613];
                
                r_data[10615] <= r_data[10614];
                
                r_data[10616] <= r_data[10615];
                
                r_data[10617] <= r_data[10616];
                
                r_data[10618] <= r_data[10617];
                
                r_data[10619] <= r_data[10618];
                
                r_data[10620] <= r_data[10619];
                
                r_data[10621] <= r_data[10620];
                
                r_data[10622] <= r_data[10621];
                
                r_data[10623] <= r_data[10622];
                
                r_data[10624] <= r_data[10623];
                
                r_data[10625] <= r_data[10624];
                
                r_data[10626] <= r_data[10625];
                
                r_data[10627] <= r_data[10626];
                
                r_data[10628] <= r_data[10627];
                
                r_data[10629] <= r_data[10628];
                
                r_data[10630] <= r_data[10629];
                
                r_data[10631] <= r_data[10630];
                
                r_data[10632] <= r_data[10631];
                
                r_data[10633] <= r_data[10632];
                
                r_data[10634] <= r_data[10633];
                
                r_data[10635] <= r_data[10634];
                
                r_data[10636] <= r_data[10635];
                
                r_data[10637] <= r_data[10636];
                
                r_data[10638] <= r_data[10637];
                
                r_data[10639] <= r_data[10638];
                
                r_data[10640] <= r_data[10639];
                
                r_data[10641] <= r_data[10640];
                
                r_data[10642] <= r_data[10641];
                
                r_data[10643] <= r_data[10642];
                
                r_data[10644] <= r_data[10643];
                
                r_data[10645] <= r_data[10644];
                
                r_data[10646] <= r_data[10645];
                
                r_data[10647] <= r_data[10646];
                
                r_data[10648] <= r_data[10647];
                
                r_data[10649] <= r_data[10648];
                
                r_data[10650] <= r_data[10649];
                
                r_data[10651] <= r_data[10650];
                
                r_data[10652] <= r_data[10651];
                
                r_data[10653] <= r_data[10652];
                
                r_data[10654] <= r_data[10653];
                
                r_data[10655] <= r_data[10654];
                
                r_data[10656] <= r_data[10655];
                
                r_data[10657] <= r_data[10656];
                
                r_data[10658] <= r_data[10657];
                
                r_data[10659] <= r_data[10658];
                
                r_data[10660] <= r_data[10659];
                
                r_data[10661] <= r_data[10660];
                
                r_data[10662] <= r_data[10661];
                
                r_data[10663] <= r_data[10662];
                
                r_data[10664] <= r_data[10663];
                
                r_data[10665] <= r_data[10664];
                
                r_data[10666] <= r_data[10665];
                
                r_data[10667] <= r_data[10666];
                
                r_data[10668] <= r_data[10667];
                
                r_data[10669] <= r_data[10668];
                
                r_data[10670] <= r_data[10669];
                
                r_data[10671] <= r_data[10670];
                
                r_data[10672] <= r_data[10671];
                
                r_data[10673] <= r_data[10672];
                
                r_data[10674] <= r_data[10673];
                
                r_data[10675] <= r_data[10674];
                
                r_data[10676] <= r_data[10675];
                
                r_data[10677] <= r_data[10676];
                
                r_data[10678] <= r_data[10677];
                
                r_data[10679] <= r_data[10678];
                
                r_data[10680] <= r_data[10679];
                
                r_data[10681] <= r_data[10680];
                
                r_data[10682] <= r_data[10681];
                
                r_data[10683] <= r_data[10682];
                
                r_data[10684] <= r_data[10683];
                
                r_data[10685] <= r_data[10684];
                
                r_data[10686] <= r_data[10685];
                
                r_data[10687] <= r_data[10686];
                
                r_data[10688] <= r_data[10687];
                
                r_data[10689] <= r_data[10688];
                
                r_data[10690] <= r_data[10689];
                
                r_data[10691] <= r_data[10690];
                
                r_data[10692] <= r_data[10691];
                
                r_data[10693] <= r_data[10692];
                
                r_data[10694] <= r_data[10693];
                
                r_data[10695] <= r_data[10694];
                
                r_data[10696] <= r_data[10695];
                
                r_data[10697] <= r_data[10696];
                
                r_data[10698] <= r_data[10697];
                
                r_data[10699] <= r_data[10698];
                
                r_data[10700] <= r_data[10699];
                
                r_data[10701] <= r_data[10700];
                
                r_data[10702] <= r_data[10701];
                
                r_data[10703] <= r_data[10702];
                
                r_data[10704] <= r_data[10703];
                
                r_data[10705] <= r_data[10704];
                
                r_data[10706] <= r_data[10705];
                
                r_data[10707] <= r_data[10706];
                
                r_data[10708] <= r_data[10707];
                
                r_data[10709] <= r_data[10708];
                
                r_data[10710] <= r_data[10709];
                
                r_data[10711] <= r_data[10710];
                
                r_data[10712] <= r_data[10711];
                
                r_data[10713] <= r_data[10712];
                
                r_data[10714] <= r_data[10713];
                
                r_data[10715] <= r_data[10714];
                
                r_data[10716] <= r_data[10715];
                
                r_data[10717] <= r_data[10716];
                
                r_data[10718] <= r_data[10717];
                
                r_data[10719] <= r_data[10718];
                
                r_data[10720] <= r_data[10719];
                
                r_data[10721] <= r_data[10720];
                
                r_data[10722] <= r_data[10721];
                
                r_data[10723] <= r_data[10722];
                
                r_data[10724] <= r_data[10723];
                
                r_data[10725] <= r_data[10724];
                
                r_data[10726] <= r_data[10725];
                
                r_data[10727] <= r_data[10726];
                
                r_data[10728] <= r_data[10727];
                
                r_data[10729] <= r_data[10728];
                
                r_data[10730] <= r_data[10729];
                
                r_data[10731] <= r_data[10730];
                
                r_data[10732] <= r_data[10731];
                
                r_data[10733] <= r_data[10732];
                
                r_data[10734] <= r_data[10733];
                
                r_data[10735] <= r_data[10734];
                
                r_data[10736] <= r_data[10735];
                
                r_data[10737] <= r_data[10736];
                
                r_data[10738] <= r_data[10737];
                
                r_data[10739] <= r_data[10738];
                
                r_data[10740] <= r_data[10739];
                
                r_data[10741] <= r_data[10740];
                
                r_data[10742] <= r_data[10741];
                
                r_data[10743] <= r_data[10742];
                
                r_data[10744] <= r_data[10743];
                
                r_data[10745] <= r_data[10744];
                
                r_data[10746] <= r_data[10745];
                
                r_data[10747] <= r_data[10746];
                
                r_data[10748] <= r_data[10747];
                
                r_data[10749] <= r_data[10748];
                
                r_data[10750] <= r_data[10749];
                
                r_data[10751] <= r_data[10750];
                
                r_data[10752] <= r_data[10751];
                
                r_data[10753] <= r_data[10752];
                
                r_data[10754] <= r_data[10753];
                
                r_data[10755] <= r_data[10754];
                
                r_data[10756] <= r_data[10755];
                
                r_data[10757] <= r_data[10756];
                
                r_data[10758] <= r_data[10757];
                
                r_data[10759] <= r_data[10758];
                
                r_data[10760] <= r_data[10759];
                
                r_data[10761] <= r_data[10760];
                
                r_data[10762] <= r_data[10761];
                
                r_data[10763] <= r_data[10762];
                
                r_data[10764] <= r_data[10763];
                
                r_data[10765] <= r_data[10764];
                
                r_data[10766] <= r_data[10765];
                
                r_data[10767] <= r_data[10766];
                
                r_data[10768] <= r_data[10767];
                
                r_data[10769] <= r_data[10768];
                
                r_data[10770] <= r_data[10769];
                
                r_data[10771] <= r_data[10770];
                
                r_data[10772] <= r_data[10771];
                
                r_data[10773] <= r_data[10772];
                
                r_data[10774] <= r_data[10773];
                
                r_data[10775] <= r_data[10774];
                
                r_data[10776] <= r_data[10775];
                
                r_data[10777] <= r_data[10776];
                
                r_data[10778] <= r_data[10777];
                
                r_data[10779] <= r_data[10778];
                
                r_data[10780] <= r_data[10779];
                
                r_data[10781] <= r_data[10780];
                
                r_data[10782] <= r_data[10781];
                
                r_data[10783] <= r_data[10782];
                
                r_data[10784] <= r_data[10783];
                
                r_data[10785] <= r_data[10784];
                
                r_data[10786] <= r_data[10785];
                
                r_data[10787] <= r_data[10786];
                
                r_data[10788] <= r_data[10787];
                
                r_data[10789] <= r_data[10788];
                
                r_data[10790] <= r_data[10789];
                
                r_data[10791] <= r_data[10790];
                
                r_data[10792] <= r_data[10791];
                
                r_data[10793] <= r_data[10792];
                
                r_data[10794] <= r_data[10793];
                
                r_data[10795] <= r_data[10794];
                
                r_data[10796] <= r_data[10795];
                
                r_data[10797] <= r_data[10796];
                
                r_data[10798] <= r_data[10797];
                
                r_data[10799] <= r_data[10798];
                
                r_data[10800] <= r_data[10799];
                
                r_data[10801] <= r_data[10800];
                
                r_data[10802] <= r_data[10801];
                
                r_data[10803] <= r_data[10802];
                
                r_data[10804] <= r_data[10803];
                
                r_data[10805] <= r_data[10804];
                
                r_data[10806] <= r_data[10805];
                
                r_data[10807] <= r_data[10806];
                
                r_data[10808] <= r_data[10807];
                
                r_data[10809] <= r_data[10808];
                
                r_data[10810] <= r_data[10809];
                
                r_data[10811] <= r_data[10810];
                
                r_data[10812] <= r_data[10811];
                
                r_data[10813] <= r_data[10812];
                
                r_data[10814] <= r_data[10813];
                
                r_data[10815] <= r_data[10814];
                
                r_data[10816] <= r_data[10815];
                
                r_data[10817] <= r_data[10816];
                
                r_data[10818] <= r_data[10817];
                
                r_data[10819] <= r_data[10818];
                
                r_data[10820] <= r_data[10819];
                
                r_data[10821] <= r_data[10820];
                
                r_data[10822] <= r_data[10821];
                
                r_data[10823] <= r_data[10822];
                
                r_data[10824] <= r_data[10823];
                
                r_data[10825] <= r_data[10824];
                
                r_data[10826] <= r_data[10825];
                
                r_data[10827] <= r_data[10826];
                
                r_data[10828] <= r_data[10827];
                
                r_data[10829] <= r_data[10828];
                
                r_data[10830] <= r_data[10829];
                
                r_data[10831] <= r_data[10830];
                
                r_data[10832] <= r_data[10831];
                
                r_data[10833] <= r_data[10832];
                
                r_data[10834] <= r_data[10833];
                
                r_data[10835] <= r_data[10834];
                
                r_data[10836] <= r_data[10835];
                
                r_data[10837] <= r_data[10836];
                
                r_data[10838] <= r_data[10837];
                
                r_data[10839] <= r_data[10838];
                
                r_data[10840] <= r_data[10839];
                
                r_data[10841] <= r_data[10840];
                
                r_data[10842] <= r_data[10841];
                
                r_data[10843] <= r_data[10842];
                
                r_data[10844] <= r_data[10843];
                
                r_data[10845] <= r_data[10844];
                
                r_data[10846] <= r_data[10845];
                
                r_data[10847] <= r_data[10846];
                
                r_data[10848] <= r_data[10847];
                
                r_data[10849] <= r_data[10848];
                
                r_data[10850] <= r_data[10849];
                
                r_data[10851] <= r_data[10850];
                
                r_data[10852] <= r_data[10851];
                
                r_data[10853] <= r_data[10852];
                
                r_data[10854] <= r_data[10853];
                
                r_data[10855] <= r_data[10854];
                
                r_data[10856] <= r_data[10855];
                
                r_data[10857] <= r_data[10856];
                
                r_data[10858] <= r_data[10857];
                
                r_data[10859] <= r_data[10858];
                
                r_data[10860] <= r_data[10859];
                
                r_data[10861] <= r_data[10860];
                
                r_data[10862] <= r_data[10861];
                
                r_data[10863] <= r_data[10862];
                
                r_data[10864] <= r_data[10863];
                
                r_data[10865] <= r_data[10864];
                
                r_data[10866] <= r_data[10865];
                
                r_data[10867] <= r_data[10866];
                
                r_data[10868] <= r_data[10867];
                
                r_data[10869] <= r_data[10868];
                
                r_data[10870] <= r_data[10869];
                
                r_data[10871] <= r_data[10870];
                
                r_data[10872] <= r_data[10871];
                
                r_data[10873] <= r_data[10872];
                
                r_data[10874] <= r_data[10873];
                
                r_data[10875] <= r_data[10874];
                
                r_data[10876] <= r_data[10875];
                
                r_data[10877] <= r_data[10876];
                
                r_data[10878] <= r_data[10877];
                
                r_data[10879] <= r_data[10878];
                
                r_data[10880] <= r_data[10879];
                
                r_data[10881] <= r_data[10880];
                
                r_data[10882] <= r_data[10881];
                
                r_data[10883] <= r_data[10882];
                
                r_data[10884] <= r_data[10883];
                
                r_data[10885] <= r_data[10884];
                
                r_data[10886] <= r_data[10885];
                
                r_data[10887] <= r_data[10886];
                
                r_data[10888] <= r_data[10887];
                
                r_data[10889] <= r_data[10888];
                
                r_data[10890] <= r_data[10889];
                
                r_data[10891] <= r_data[10890];
                
                r_data[10892] <= r_data[10891];
                
                r_data[10893] <= r_data[10892];
                
                r_data[10894] <= r_data[10893];
                
                r_data[10895] <= r_data[10894];
                
                r_data[10896] <= r_data[10895];
                
                r_data[10897] <= r_data[10896];
                
                r_data[10898] <= r_data[10897];
                
                r_data[10899] <= r_data[10898];
                
                r_data[10900] <= r_data[10899];
                
                r_data[10901] <= r_data[10900];
                
                r_data[10902] <= r_data[10901];
                
                r_data[10903] <= r_data[10902];
                
                r_data[10904] <= r_data[10903];
                
                r_data[10905] <= r_data[10904];
                
                r_data[10906] <= r_data[10905];
                
                r_data[10907] <= r_data[10906];
                
                r_data[10908] <= r_data[10907];
                
                r_data[10909] <= r_data[10908];
                
                r_data[10910] <= r_data[10909];
                
                r_data[10911] <= r_data[10910];
                
                r_data[10912] <= r_data[10911];
                
                r_data[10913] <= r_data[10912];
                
                r_data[10914] <= r_data[10913];
                
                r_data[10915] <= r_data[10914];
                
                r_data[10916] <= r_data[10915];
                
                r_data[10917] <= r_data[10916];
                
                r_data[10918] <= r_data[10917];
                
                r_data[10919] <= r_data[10918];
                
                r_data[10920] <= r_data[10919];
                
                r_data[10921] <= r_data[10920];
                
                r_data[10922] <= r_data[10921];
                
                r_data[10923] <= r_data[10922];
                
                r_data[10924] <= r_data[10923];
                
                r_data[10925] <= r_data[10924];
                
                r_data[10926] <= r_data[10925];
                
                r_data[10927] <= r_data[10926];
                
                r_data[10928] <= r_data[10927];
                
                r_data[10929] <= r_data[10928];
                
                r_data[10930] <= r_data[10929];
                
                r_data[10931] <= r_data[10930];
                
                r_data[10932] <= r_data[10931];
                
                r_data[10933] <= r_data[10932];
                
                r_data[10934] <= r_data[10933];
                
                r_data[10935] <= r_data[10934];
                
                r_data[10936] <= r_data[10935];
                
                r_data[10937] <= r_data[10936];
                
                r_data[10938] <= r_data[10937];
                
                r_data[10939] <= r_data[10938];
                
                r_data[10940] <= r_data[10939];
                
                r_data[10941] <= r_data[10940];
                
                r_data[10942] <= r_data[10941];
                
                r_data[10943] <= r_data[10942];
                
                r_data[10944] <= r_data[10943];
                
                r_data[10945] <= r_data[10944];
                
                r_data[10946] <= r_data[10945];
                
                r_data[10947] <= r_data[10946];
                
                r_data[10948] <= r_data[10947];
                
                r_data[10949] <= r_data[10948];
                
                r_data[10950] <= r_data[10949];
                
                r_data[10951] <= r_data[10950];
                
                r_data[10952] <= r_data[10951];
                
                r_data[10953] <= r_data[10952];
                
                r_data[10954] <= r_data[10953];
                
                r_data[10955] <= r_data[10954];
                
                r_data[10956] <= r_data[10955];
                
                r_data[10957] <= r_data[10956];
                
                r_data[10958] <= r_data[10957];
                
                r_data[10959] <= r_data[10958];
                
                r_data[10960] <= r_data[10959];
                
                r_data[10961] <= r_data[10960];
                
                r_data[10962] <= r_data[10961];
                
                r_data[10963] <= r_data[10962];
                
                r_data[10964] <= r_data[10963];
                
                r_data[10965] <= r_data[10964];
                
                r_data[10966] <= r_data[10965];
                
                r_data[10967] <= r_data[10966];
                
                r_data[10968] <= r_data[10967];
                
                r_data[10969] <= r_data[10968];
                
                r_data[10970] <= r_data[10969];
                
                r_data[10971] <= r_data[10970];
                
                r_data[10972] <= r_data[10971];
                
                r_data[10973] <= r_data[10972];
                
                r_data[10974] <= r_data[10973];
                
                r_data[10975] <= r_data[10974];
                
                r_data[10976] <= r_data[10975];
                
                r_data[10977] <= r_data[10976];
                
                r_data[10978] <= r_data[10977];
                
                r_data[10979] <= r_data[10978];
                
                r_data[10980] <= r_data[10979];
                
                r_data[10981] <= r_data[10980];
                
                r_data[10982] <= r_data[10981];
                
                r_data[10983] <= r_data[10982];
                
                r_data[10984] <= r_data[10983];
                
                r_data[10985] <= r_data[10984];
                
                r_data[10986] <= r_data[10985];
                
                r_data[10987] <= r_data[10986];
                
                r_data[10988] <= r_data[10987];
                
                r_data[10989] <= r_data[10988];
                
                r_data[10990] <= r_data[10989];
                
                r_data[10991] <= r_data[10990];
                
                r_data[10992] <= r_data[10991];
                
                r_data[10993] <= r_data[10992];
                
                r_data[10994] <= r_data[10993];
                
                r_data[10995] <= r_data[10994];
                
                r_data[10996] <= r_data[10995];
                
                r_data[10997] <= r_data[10996];
                
                r_data[10998] <= r_data[10997];
                
                r_data[10999] <= r_data[10998];
                
                r_data[11000] <= r_data[10999];
                
                r_data[11001] <= r_data[11000];
                
                r_data[11002] <= r_data[11001];
                
                r_data[11003] <= r_data[11002];
                
                r_data[11004] <= r_data[11003];
                
                r_data[11005] <= r_data[11004];
                
                r_data[11006] <= r_data[11005];
                
                r_data[11007] <= r_data[11006];
                
                r_data[11008] <= r_data[11007];
                
                r_data[11009] <= r_data[11008];
                
                r_data[11010] <= r_data[11009];
                
                r_data[11011] <= r_data[11010];
                
                r_data[11012] <= r_data[11011];
                
                r_data[11013] <= r_data[11012];
                
                r_data[11014] <= r_data[11013];
                
                r_data[11015] <= r_data[11014];
                
                r_data[11016] <= r_data[11015];
                
                r_data[11017] <= r_data[11016];
                
                r_data[11018] <= r_data[11017];
                
                r_data[11019] <= r_data[11018];
                
                r_data[11020] <= r_data[11019];
                
                r_data[11021] <= r_data[11020];
                
                r_data[11022] <= r_data[11021];
                
                r_data[11023] <= r_data[11022];
                
                r_data[11024] <= r_data[11023];
                
                r_data[11025] <= r_data[11024];
                
                r_data[11026] <= r_data[11025];
                
                r_data[11027] <= r_data[11026];
                
                r_data[11028] <= r_data[11027];
                
                r_data[11029] <= r_data[11028];
                
                r_data[11030] <= r_data[11029];
                
                r_data[11031] <= r_data[11030];
                
                r_data[11032] <= r_data[11031];
                
                r_data[11033] <= r_data[11032];
                
                r_data[11034] <= r_data[11033];
                
                r_data[11035] <= r_data[11034];
                
                r_data[11036] <= r_data[11035];
                
                r_data[11037] <= r_data[11036];
                
                r_data[11038] <= r_data[11037];
                
                r_data[11039] <= r_data[11038];
                
                r_data[11040] <= r_data[11039];
                
                r_data[11041] <= r_data[11040];
                
                r_data[11042] <= r_data[11041];
                
                r_data[11043] <= r_data[11042];
                
                r_data[11044] <= r_data[11043];
                
                r_data[11045] <= r_data[11044];
                
                r_data[11046] <= r_data[11045];
                
                r_data[11047] <= r_data[11046];
                
                r_data[11048] <= r_data[11047];
                
                r_data[11049] <= r_data[11048];
                
                r_data[11050] <= r_data[11049];
                
                r_data[11051] <= r_data[11050];
                
                r_data[11052] <= r_data[11051];
                
                r_data[11053] <= r_data[11052];
                
                r_data[11054] <= r_data[11053];
                
                r_data[11055] <= r_data[11054];
                
                r_data[11056] <= r_data[11055];
                
                r_data[11057] <= r_data[11056];
                
                r_data[11058] <= r_data[11057];
                
                r_data[11059] <= r_data[11058];
                
                r_data[11060] <= r_data[11059];
                
                r_data[11061] <= r_data[11060];
                
                r_data[11062] <= r_data[11061];
                
                r_data[11063] <= r_data[11062];
                
                r_data[11064] <= r_data[11063];
                
                r_data[11065] <= r_data[11064];
                
                r_data[11066] <= r_data[11065];
                
                r_data[11067] <= r_data[11066];
                
                r_data[11068] <= r_data[11067];
                
                r_data[11069] <= r_data[11068];
                
                r_data[11070] <= r_data[11069];
                
                r_data[11071] <= r_data[11070];
                
                r_data[11072] <= r_data[11071];
                
                r_data[11073] <= r_data[11072];
                
                r_data[11074] <= r_data[11073];
                
                r_data[11075] <= r_data[11074];
                
                r_data[11076] <= r_data[11075];
                
                r_data[11077] <= r_data[11076];
                
                r_data[11078] <= r_data[11077];
                
                r_data[11079] <= r_data[11078];
                
                r_data[11080] <= r_data[11079];
                
                r_data[11081] <= r_data[11080];
                
                r_data[11082] <= r_data[11081];
                
                r_data[11083] <= r_data[11082];
                
                r_data[11084] <= r_data[11083];
                
                r_data[11085] <= r_data[11084];
                
                r_data[11086] <= r_data[11085];
                
                r_data[11087] <= r_data[11086];
                
                r_data[11088] <= r_data[11087];
                
                r_data[11089] <= r_data[11088];
                
                r_data[11090] <= r_data[11089];
                
                r_data[11091] <= r_data[11090];
                
                r_data[11092] <= r_data[11091];
                
                r_data[11093] <= r_data[11092];
                
                r_data[11094] <= r_data[11093];
                
                r_data[11095] <= r_data[11094];
                
                r_data[11096] <= r_data[11095];
                
                r_data[11097] <= r_data[11096];
                
                r_data[11098] <= r_data[11097];
                
                r_data[11099] <= r_data[11098];
                
                r_data[11100] <= r_data[11099];
                
                r_data[11101] <= r_data[11100];
                
                r_data[11102] <= r_data[11101];
                
                r_data[11103] <= r_data[11102];
                
                r_data[11104] <= r_data[11103];
                
                r_data[11105] <= r_data[11104];
                
                r_data[11106] <= r_data[11105];
                
                r_data[11107] <= r_data[11106];
                
                r_data[11108] <= r_data[11107];
                
                r_data[11109] <= r_data[11108];
                
                r_data[11110] <= r_data[11109];
                
                r_data[11111] <= r_data[11110];
                
                r_data[11112] <= r_data[11111];
                
                r_data[11113] <= r_data[11112];
                
                r_data[11114] <= r_data[11113];
                
                r_data[11115] <= r_data[11114];
                
                r_data[11116] <= r_data[11115];
                
                r_data[11117] <= r_data[11116];
                
                r_data[11118] <= r_data[11117];
                
                r_data[11119] <= r_data[11118];
                
                r_data[11120] <= r_data[11119];
                
                r_data[11121] <= r_data[11120];
                
                r_data[11122] <= r_data[11121];
                
                r_data[11123] <= r_data[11122];
                
                r_data[11124] <= r_data[11123];
                
                r_data[11125] <= r_data[11124];
                
                r_data[11126] <= r_data[11125];
                
                r_data[11127] <= r_data[11126];
                
                r_data[11128] <= r_data[11127];
                
                r_data[11129] <= r_data[11128];
                
                r_data[11130] <= r_data[11129];
                
                r_data[11131] <= r_data[11130];
                
                r_data[11132] <= r_data[11131];
                
                r_data[11133] <= r_data[11132];
                
                r_data[11134] <= r_data[11133];
                
                r_data[11135] <= r_data[11134];
                
                r_data[11136] <= r_data[11135];
                
                r_data[11137] <= r_data[11136];
                
                r_data[11138] <= r_data[11137];
                
                r_data[11139] <= r_data[11138];
                
                r_data[11140] <= r_data[11139];
                
                r_data[11141] <= r_data[11140];
                
                r_data[11142] <= r_data[11141];
                
                r_data[11143] <= r_data[11142];
                
                r_data[11144] <= r_data[11143];
                
                r_data[11145] <= r_data[11144];
                
                r_data[11146] <= r_data[11145];
                
                r_data[11147] <= r_data[11146];
                
                r_data[11148] <= r_data[11147];
                
                r_data[11149] <= r_data[11148];
                
                r_data[11150] <= r_data[11149];
                
                r_data[11151] <= r_data[11150];
                
                r_data[11152] <= r_data[11151];
                
                r_data[11153] <= r_data[11152];
                
                r_data[11154] <= r_data[11153];
                
                r_data[11155] <= r_data[11154];
                
                r_data[11156] <= r_data[11155];
                
                r_data[11157] <= r_data[11156];
                
                r_data[11158] <= r_data[11157];
                
                r_data[11159] <= r_data[11158];
                
                r_data[11160] <= r_data[11159];
                
                r_data[11161] <= r_data[11160];
                
                r_data[11162] <= r_data[11161];
                
                r_data[11163] <= r_data[11162];
                
                r_data[11164] <= r_data[11163];
                
                r_data[11165] <= r_data[11164];
                
                r_data[11166] <= r_data[11165];
                
                r_data[11167] <= r_data[11166];
                
                r_data[11168] <= r_data[11167];
                
                r_data[11169] <= r_data[11168];
                
                r_data[11170] <= r_data[11169];
                
                r_data[11171] <= r_data[11170];
                
                r_data[11172] <= r_data[11171];
                
                r_data[11173] <= r_data[11172];
                
                r_data[11174] <= r_data[11173];
                
                r_data[11175] <= r_data[11174];
                
                r_data[11176] <= r_data[11175];
                
                r_data[11177] <= r_data[11176];
                
                r_data[11178] <= r_data[11177];
                
                r_data[11179] <= r_data[11178];
                
                r_data[11180] <= r_data[11179];
                
                r_data[11181] <= r_data[11180];
                
                r_data[11182] <= r_data[11181];
                
                r_data[11183] <= r_data[11182];
                
                r_data[11184] <= r_data[11183];
                
                r_data[11185] <= r_data[11184];
                
                r_data[11186] <= r_data[11185];
                
                r_data[11187] <= r_data[11186];
                
                r_data[11188] <= r_data[11187];
                
                r_data[11189] <= r_data[11188];
                
                r_data[11190] <= r_data[11189];
                
                r_data[11191] <= r_data[11190];
                
                r_data[11192] <= r_data[11191];
                
                r_data[11193] <= r_data[11192];
                
                r_data[11194] <= r_data[11193];
                
                r_data[11195] <= r_data[11194];
                
                r_data[11196] <= r_data[11195];
                
                r_data[11197] <= r_data[11196];
                
                r_data[11198] <= r_data[11197];
                
                r_data[11199] <= r_data[11198];
                
                r_data[11200] <= r_data[11199];
                
                r_data[11201] <= r_data[11200];
                
                r_data[11202] <= r_data[11201];
                
                r_data[11203] <= r_data[11202];
                
                r_data[11204] <= r_data[11203];
                
                r_data[11205] <= r_data[11204];
                
                r_data[11206] <= r_data[11205];
                
                r_data[11207] <= r_data[11206];
                
                r_data[11208] <= r_data[11207];
                
                r_data[11209] <= r_data[11208];
                
                r_data[11210] <= r_data[11209];
                
                r_data[11211] <= r_data[11210];
                
                r_data[11212] <= r_data[11211];
                
                r_data[11213] <= r_data[11212];
                
                r_data[11214] <= r_data[11213];
                
                r_data[11215] <= r_data[11214];
                
                r_data[11216] <= r_data[11215];
                
                r_data[11217] <= r_data[11216];
                
                r_data[11218] <= r_data[11217];
                
                r_data[11219] <= r_data[11218];
                
                r_data[11220] <= r_data[11219];
                
                r_data[11221] <= r_data[11220];
                
                r_data[11222] <= r_data[11221];
                
                r_data[11223] <= r_data[11222];
                
                r_data[11224] <= r_data[11223];
                
                r_data[11225] <= r_data[11224];
                
                r_data[11226] <= r_data[11225];
                
                r_data[11227] <= r_data[11226];
                
                r_data[11228] <= r_data[11227];
                
                r_data[11229] <= r_data[11228];
                
                r_data[11230] <= r_data[11229];
                
                r_data[11231] <= r_data[11230];
                
                r_data[11232] <= r_data[11231];
                
                r_data[11233] <= r_data[11232];
                
                r_data[11234] <= r_data[11233];
                
                r_data[11235] <= r_data[11234];
                
                r_data[11236] <= r_data[11235];
                
                r_data[11237] <= r_data[11236];
                
                r_data[11238] <= r_data[11237];
                
                r_data[11239] <= r_data[11238];
                
                r_data[11240] <= r_data[11239];
                
                r_data[11241] <= r_data[11240];
                
                r_data[11242] <= r_data[11241];
                
                r_data[11243] <= r_data[11242];
                
                r_data[11244] <= r_data[11243];
                
                r_data[11245] <= r_data[11244];
                
                r_data[11246] <= r_data[11245];
                
                r_data[11247] <= r_data[11246];
                
                r_data[11248] <= r_data[11247];
                
                r_data[11249] <= r_data[11248];
                
                r_data[11250] <= r_data[11249];
                
                r_data[11251] <= r_data[11250];
                
                r_data[11252] <= r_data[11251];
                
                r_data[11253] <= r_data[11252];
                
                r_data[11254] <= r_data[11253];
                
                r_data[11255] <= r_data[11254];
                
                r_data[11256] <= r_data[11255];
                
                r_data[11257] <= r_data[11256];
                
                r_data[11258] <= r_data[11257];
                
                r_data[11259] <= r_data[11258];
                
                r_data[11260] <= r_data[11259];
                
                r_data[11261] <= r_data[11260];
                
                r_data[11262] <= r_data[11261];
                
                r_data[11263] <= r_data[11262];
                
                r_data[11264] <= r_data[11263];
                
                r_data[11265] <= r_data[11264];
                
                r_data[11266] <= r_data[11265];
                
                r_data[11267] <= r_data[11266];
                
                r_data[11268] <= r_data[11267];
                
                r_data[11269] <= r_data[11268];
                
                r_data[11270] <= r_data[11269];
                
                r_data[11271] <= r_data[11270];
                
                r_data[11272] <= r_data[11271];
                
                r_data[11273] <= r_data[11272];
                
                r_data[11274] <= r_data[11273];
                
                r_data[11275] <= r_data[11274];
                
                r_data[11276] <= r_data[11275];
                
                r_data[11277] <= r_data[11276];
                
                r_data[11278] <= r_data[11277];
                
                r_data[11279] <= r_data[11278];
                
                r_data[11280] <= r_data[11279];
                
                r_data[11281] <= r_data[11280];
                
                r_data[11282] <= r_data[11281];
                
                r_data[11283] <= r_data[11282];
                
                r_data[11284] <= r_data[11283];
                
                r_data[11285] <= r_data[11284];
                
                r_data[11286] <= r_data[11285];
                
                r_data[11287] <= r_data[11286];
                
                r_data[11288] <= r_data[11287];
                
                r_data[11289] <= r_data[11288];
                
                r_data[11290] <= r_data[11289];
                
                r_data[11291] <= r_data[11290];
                
                r_data[11292] <= r_data[11291];
                
                r_data[11293] <= r_data[11292];
                
                r_data[11294] <= r_data[11293];
                
                r_data[11295] <= r_data[11294];
                
                r_data[11296] <= r_data[11295];
                
                r_data[11297] <= r_data[11296];
                
                r_data[11298] <= r_data[11297];
                
                r_data[11299] <= r_data[11298];
                
                r_data[11300] <= r_data[11299];
                
                r_data[11301] <= r_data[11300];
                
                r_data[11302] <= r_data[11301];
                
                r_data[11303] <= r_data[11302];
                
                r_data[11304] <= r_data[11303];
                
                r_data[11305] <= r_data[11304];
                
                r_data[11306] <= r_data[11305];
                
                r_data[11307] <= r_data[11306];
                
                r_data[11308] <= r_data[11307];
                
                r_data[11309] <= r_data[11308];
                
                r_data[11310] <= r_data[11309];
                
                r_data[11311] <= r_data[11310];
                
                r_data[11312] <= r_data[11311];
                
                r_data[11313] <= r_data[11312];
                
                r_data[11314] <= r_data[11313];
                
                r_data[11315] <= r_data[11314];
                
                r_data[11316] <= r_data[11315];
                
                r_data[11317] <= r_data[11316];
                
                r_data[11318] <= r_data[11317];
                
                r_data[11319] <= r_data[11318];
                
                r_data[11320] <= r_data[11319];
                
                r_data[11321] <= r_data[11320];
                
                r_data[11322] <= r_data[11321];
                
                r_data[11323] <= r_data[11322];
                
                r_data[11324] <= r_data[11323];
                
                r_data[11325] <= r_data[11324];
                
                r_data[11326] <= r_data[11325];
                
                r_data[11327] <= r_data[11326];
                
                r_data[11328] <= r_data[11327];
                
                r_data[11329] <= r_data[11328];
                
                r_data[11330] <= r_data[11329];
                
                r_data[11331] <= r_data[11330];
                
                r_data[11332] <= r_data[11331];
                
                r_data[11333] <= r_data[11332];
                
                r_data[11334] <= r_data[11333];
                
                r_data[11335] <= r_data[11334];
                
                r_data[11336] <= r_data[11335];
                
                r_data[11337] <= r_data[11336];
                
                r_data[11338] <= r_data[11337];
                
                r_data[11339] <= r_data[11338];
                
                r_data[11340] <= r_data[11339];
                
                r_data[11341] <= r_data[11340];
                
                r_data[11342] <= r_data[11341];
                
                r_data[11343] <= r_data[11342];
                
                r_data[11344] <= r_data[11343];
                
                r_data[11345] <= r_data[11344];
                
                r_data[11346] <= r_data[11345];
                
                r_data[11347] <= r_data[11346];
                
                r_data[11348] <= r_data[11347];
                
                r_data[11349] <= r_data[11348];
                
                r_data[11350] <= r_data[11349];
                
                r_data[11351] <= r_data[11350];
                
                r_data[11352] <= r_data[11351];
                
                r_data[11353] <= r_data[11352];
                
                r_data[11354] <= r_data[11353];
                
                r_data[11355] <= r_data[11354];
                
                r_data[11356] <= r_data[11355];
                
                r_data[11357] <= r_data[11356];
                
                r_data[11358] <= r_data[11357];
                
                r_data[11359] <= r_data[11358];
                
                r_data[11360] <= r_data[11359];
                
                r_data[11361] <= r_data[11360];
                
                r_data[11362] <= r_data[11361];
                
                r_data[11363] <= r_data[11362];
                
                r_data[11364] <= r_data[11363];
                
                r_data[11365] <= r_data[11364];
                
                r_data[11366] <= r_data[11365];
                
                r_data[11367] <= r_data[11366];
                
                r_data[11368] <= r_data[11367];
                
                r_data[11369] <= r_data[11368];
                
                r_data[11370] <= r_data[11369];
                
                r_data[11371] <= r_data[11370];
                
                r_data[11372] <= r_data[11371];
                
                r_data[11373] <= r_data[11372];
                
                r_data[11374] <= r_data[11373];
                
                r_data[11375] <= r_data[11374];
                
                r_data[11376] <= r_data[11375];
                
                r_data[11377] <= r_data[11376];
                
                r_data[11378] <= r_data[11377];
                
                r_data[11379] <= r_data[11378];
                
                r_data[11380] <= r_data[11379];
                
                r_data[11381] <= r_data[11380];
                
                r_data[11382] <= r_data[11381];
                
                r_data[11383] <= r_data[11382];
                
                r_data[11384] <= r_data[11383];
                
                r_data[11385] <= r_data[11384];
                
                r_data[11386] <= r_data[11385];
                
                r_data[11387] <= r_data[11386];
                
                r_data[11388] <= r_data[11387];
                
                r_data[11389] <= r_data[11388];
                
                r_data[11390] <= r_data[11389];
                
                r_data[11391] <= r_data[11390];
                
                r_data[11392] <= r_data[11391];
                
                r_data[11393] <= r_data[11392];
                
                r_data[11394] <= r_data[11393];
                
                r_data[11395] <= r_data[11394];
                
                r_data[11396] <= r_data[11395];
                
                r_data[11397] <= r_data[11396];
                
                r_data[11398] <= r_data[11397];
                
                r_data[11399] <= r_data[11398];
                
                r_data[11400] <= r_data[11399];
                
                r_data[11401] <= r_data[11400];
                
                r_data[11402] <= r_data[11401];
                
                r_data[11403] <= r_data[11402];
                
                r_data[11404] <= r_data[11403];
                
                r_data[11405] <= r_data[11404];
                
                r_data[11406] <= r_data[11405];
                
                r_data[11407] <= r_data[11406];
                
                r_data[11408] <= r_data[11407];
                
                r_data[11409] <= r_data[11408];
                
                r_data[11410] <= r_data[11409];
                
                r_data[11411] <= r_data[11410];
                
                r_data[11412] <= r_data[11411];
                
                r_data[11413] <= r_data[11412];
                
                r_data[11414] <= r_data[11413];
                
                r_data[11415] <= r_data[11414];
                
                r_data[11416] <= r_data[11415];
                
                r_data[11417] <= r_data[11416];
                
                r_data[11418] <= r_data[11417];
                
                r_data[11419] <= r_data[11418];
                
                r_data[11420] <= r_data[11419];
                
                r_data[11421] <= r_data[11420];
                
                r_data[11422] <= r_data[11421];
                
                r_data[11423] <= r_data[11422];
                
                r_data[11424] <= r_data[11423];
                
                r_data[11425] <= r_data[11424];
                
                r_data[11426] <= r_data[11425];
                
                r_data[11427] <= r_data[11426];
                
                r_data[11428] <= r_data[11427];
                
                r_data[11429] <= r_data[11428];
                
                r_data[11430] <= r_data[11429];
                
                r_data[11431] <= r_data[11430];
                
                r_data[11432] <= r_data[11431];
                
                r_data[11433] <= r_data[11432];
                
                r_data[11434] <= r_data[11433];
                
                r_data[11435] <= r_data[11434];
                
                r_data[11436] <= r_data[11435];
                
                r_data[11437] <= r_data[11436];
                
                r_data[11438] <= r_data[11437];
                
                r_data[11439] <= r_data[11438];
                
                r_data[11440] <= r_data[11439];
                
                r_data[11441] <= r_data[11440];
                
                r_data[11442] <= r_data[11441];
                
                r_data[11443] <= r_data[11442];
                
                r_data[11444] <= r_data[11443];
                
                r_data[11445] <= r_data[11444];
                
                r_data[11446] <= r_data[11445];
                
                r_data[11447] <= r_data[11446];
                
                r_data[11448] <= r_data[11447];
                
                r_data[11449] <= r_data[11448];
                
                r_data[11450] <= r_data[11449];
                
                r_data[11451] <= r_data[11450];
                
                r_data[11452] <= r_data[11451];
                
                r_data[11453] <= r_data[11452];
                
                r_data[11454] <= r_data[11453];
                
                r_data[11455] <= r_data[11454];
                
                r_data[11456] <= r_data[11455];
                
                r_data[11457] <= r_data[11456];
                
                r_data[11458] <= r_data[11457];
                
                r_data[11459] <= r_data[11458];
                
                r_data[11460] <= r_data[11459];
                
                r_data[11461] <= r_data[11460];
                
                r_data[11462] <= r_data[11461];
                
                r_data[11463] <= r_data[11462];
                
                r_data[11464] <= r_data[11463];
                
                r_data[11465] <= r_data[11464];
                
                r_data[11466] <= r_data[11465];
                
                r_data[11467] <= r_data[11466];
                
                r_data[11468] <= r_data[11467];
                
                r_data[11469] <= r_data[11468];
                
                r_data[11470] <= r_data[11469];
                
                r_data[11471] <= r_data[11470];
                
                r_data[11472] <= r_data[11471];
                
                r_data[11473] <= r_data[11472];
                
                r_data[11474] <= r_data[11473];
                
                r_data[11475] <= r_data[11474];
                
                r_data[11476] <= r_data[11475];
                
                r_data[11477] <= r_data[11476];
                
                r_data[11478] <= r_data[11477];
                
                r_data[11479] <= r_data[11478];
                
                r_data[11480] <= r_data[11479];
                
                r_data[11481] <= r_data[11480];
                
                r_data[11482] <= r_data[11481];
                
                r_data[11483] <= r_data[11482];
                
                r_data[11484] <= r_data[11483];
                
                r_data[11485] <= r_data[11484];
                
                r_data[11486] <= r_data[11485];
                
                r_data[11487] <= r_data[11486];
                
                r_data[11488] <= r_data[11487];
                
                r_data[11489] <= r_data[11488];
                
                r_data[11490] <= r_data[11489];
                
                r_data[11491] <= r_data[11490];
                
                r_data[11492] <= r_data[11491];
                
                r_data[11493] <= r_data[11492];
                
                r_data[11494] <= r_data[11493];
                
                r_data[11495] <= r_data[11494];
                
                r_data[11496] <= r_data[11495];
                
                r_data[11497] <= r_data[11496];
                
                r_data[11498] <= r_data[11497];
                
                r_data[11499] <= r_data[11498];
                
                r_data[11500] <= r_data[11499];
                
                r_data[11501] <= r_data[11500];
                
                r_data[11502] <= r_data[11501];
                
                r_data[11503] <= r_data[11502];
                
                r_data[11504] <= r_data[11503];
                
                r_data[11505] <= r_data[11504];
                
                r_data[11506] <= r_data[11505];
                
                r_data[11507] <= r_data[11506];
                
                r_data[11508] <= r_data[11507];
                
                r_data[11509] <= r_data[11508];
                
                r_data[11510] <= r_data[11509];
                
                r_data[11511] <= r_data[11510];
                
                r_data[11512] <= r_data[11511];
                
                r_data[11513] <= r_data[11512];
                
                r_data[11514] <= r_data[11513];
                
                r_data[11515] <= r_data[11514];
                
                r_data[11516] <= r_data[11515];
                
                r_data[11517] <= r_data[11516];
                
                r_data[11518] <= r_data[11517];
                
                r_data[11519] <= r_data[11518];
                
                r_data[11520] <= r_data[11519];
                
                r_data[11521] <= r_data[11520];
                
                r_data[11522] <= r_data[11521];
                
                r_data[11523] <= r_data[11522];
                
                r_data[11524] <= r_data[11523];
                
                r_data[11525] <= r_data[11524];
                
                r_data[11526] <= r_data[11525];
                
                r_data[11527] <= r_data[11526];
                
                r_data[11528] <= r_data[11527];
                
                r_data[11529] <= r_data[11528];
                
                r_data[11530] <= r_data[11529];
                
                r_data[11531] <= r_data[11530];
                
                r_data[11532] <= r_data[11531];
                
                r_data[11533] <= r_data[11532];
                
                r_data[11534] <= r_data[11533];
                
                r_data[11535] <= r_data[11534];
                
                r_data[11536] <= r_data[11535];
                
                r_data[11537] <= r_data[11536];
                
                r_data[11538] <= r_data[11537];
                
                r_data[11539] <= r_data[11538];
                
                r_data[11540] <= r_data[11539];
                
                r_data[11541] <= r_data[11540];
                
                r_data[11542] <= r_data[11541];
                
                r_data[11543] <= r_data[11542];
                
                r_data[11544] <= r_data[11543];
                
                r_data[11545] <= r_data[11544];
                
                r_data[11546] <= r_data[11545];
                
                r_data[11547] <= r_data[11546];
                
                r_data[11548] <= r_data[11547];
                
                r_data[11549] <= r_data[11548];
                
                r_data[11550] <= r_data[11549];
                
                r_data[11551] <= r_data[11550];
                
                r_data[11552] <= r_data[11551];
                
                r_data[11553] <= r_data[11552];
                
                r_data[11554] <= r_data[11553];
                
                r_data[11555] <= r_data[11554];
                
                r_data[11556] <= r_data[11555];
                
                r_data[11557] <= r_data[11556];
                
                r_data[11558] <= r_data[11557];
                
                r_data[11559] <= r_data[11558];
                
                r_data[11560] <= r_data[11559];
                
                r_data[11561] <= r_data[11560];
                
                r_data[11562] <= r_data[11561];
                
                r_data[11563] <= r_data[11562];
                
                r_data[11564] <= r_data[11563];
                
                r_data[11565] <= r_data[11564];
                
                r_data[11566] <= r_data[11565];
                
                r_data[11567] <= r_data[11566];
                
                r_data[11568] <= r_data[11567];
                
                r_data[11569] <= r_data[11568];
                
                r_data[11570] <= r_data[11569];
                
                r_data[11571] <= r_data[11570];
                
                r_data[11572] <= r_data[11571];
                
                r_data[11573] <= r_data[11572];
                
                r_data[11574] <= r_data[11573];
                
                r_data[11575] <= r_data[11574];
                
                r_data[11576] <= r_data[11575];
                
                r_data[11577] <= r_data[11576];
                
                r_data[11578] <= r_data[11577];
                
                r_data[11579] <= r_data[11578];
                
                r_data[11580] <= r_data[11579];
                
                r_data[11581] <= r_data[11580];
                
                r_data[11582] <= r_data[11581];
                
                r_data[11583] <= r_data[11582];
                
                r_data[11584] <= r_data[11583];
                
                r_data[11585] <= r_data[11584];
                
                r_data[11586] <= r_data[11585];
                
                r_data[11587] <= r_data[11586];
                
                r_data[11588] <= r_data[11587];
                
                r_data[11589] <= r_data[11588];
                
                r_data[11590] <= r_data[11589];
                
                r_data[11591] <= r_data[11590];
                
                r_data[11592] <= r_data[11591];
                
                r_data[11593] <= r_data[11592];
                
                r_data[11594] <= r_data[11593];
                
                r_data[11595] <= r_data[11594];
                
                r_data[11596] <= r_data[11595];
                
                r_data[11597] <= r_data[11596];
                
                r_data[11598] <= r_data[11597];
                
                r_data[11599] <= r_data[11598];
                
                r_data[11600] <= r_data[11599];
                
                r_data[11601] <= r_data[11600];
                
                r_data[11602] <= r_data[11601];
                
                r_data[11603] <= r_data[11602];
                
                r_data[11604] <= r_data[11603];
                
                r_data[11605] <= r_data[11604];
                
                r_data[11606] <= r_data[11605];
                
                r_data[11607] <= r_data[11606];
                
                r_data[11608] <= r_data[11607];
                
                r_data[11609] <= r_data[11608];
                
                r_data[11610] <= r_data[11609];
                
                r_data[11611] <= r_data[11610];
                
                r_data[11612] <= r_data[11611];
                
                r_data[11613] <= r_data[11612];
                
                r_data[11614] <= r_data[11613];
                
                r_data[11615] <= r_data[11614];
                
                r_data[11616] <= r_data[11615];
                
                r_data[11617] <= r_data[11616];
                
                r_data[11618] <= r_data[11617];
                
                r_data[11619] <= r_data[11618];
                
                r_data[11620] <= r_data[11619];
                
                r_data[11621] <= r_data[11620];
                
                r_data[11622] <= r_data[11621];
                
                r_data[11623] <= r_data[11622];
                
                r_data[11624] <= r_data[11623];
                
                r_data[11625] <= r_data[11624];
                
                r_data[11626] <= r_data[11625];
                
                r_data[11627] <= r_data[11626];
                
                r_data[11628] <= r_data[11627];
                
                r_data[11629] <= r_data[11628];
                
                r_data[11630] <= r_data[11629];
                
                r_data[11631] <= r_data[11630];
                
                r_data[11632] <= r_data[11631];
                
                r_data[11633] <= r_data[11632];
                
                r_data[11634] <= r_data[11633];
                
                r_data[11635] <= r_data[11634];
                
                r_data[11636] <= r_data[11635];
                
                r_data[11637] <= r_data[11636];
                
                r_data[11638] <= r_data[11637];
                
                r_data[11639] <= r_data[11638];
                
                r_data[11640] <= r_data[11639];
                
                r_data[11641] <= r_data[11640];
                
                r_data[11642] <= r_data[11641];
                
                r_data[11643] <= r_data[11642];
                
                r_data[11644] <= r_data[11643];
                
                r_data[11645] <= r_data[11644];
                
                r_data[11646] <= r_data[11645];
                
                r_data[11647] <= r_data[11646];
                
                r_data[11648] <= r_data[11647];
                
                r_data[11649] <= r_data[11648];
                
                r_data[11650] <= r_data[11649];
                
                r_data[11651] <= r_data[11650];
                
                r_data[11652] <= r_data[11651];
                
                r_data[11653] <= r_data[11652];
                
                r_data[11654] <= r_data[11653];
                
                r_data[11655] <= r_data[11654];
                
                r_data[11656] <= r_data[11655];
                
                r_data[11657] <= r_data[11656];
                
                r_data[11658] <= r_data[11657];
                
                r_data[11659] <= r_data[11658];
                
                r_data[11660] <= r_data[11659];
                
                r_data[11661] <= r_data[11660];
                
                r_data[11662] <= r_data[11661];
                
                r_data[11663] <= r_data[11662];
                
                r_data[11664] <= r_data[11663];
                
                r_data[11665] <= r_data[11664];
                
                r_data[11666] <= r_data[11665];
                
                r_data[11667] <= r_data[11666];
                
                r_data[11668] <= r_data[11667];
                
                r_data[11669] <= r_data[11668];
                
                r_data[11670] <= r_data[11669];
                
                r_data[11671] <= r_data[11670];
                
                r_data[11672] <= r_data[11671];
                
                r_data[11673] <= r_data[11672];
                
                r_data[11674] <= r_data[11673];
                
                r_data[11675] <= r_data[11674];
                
                r_data[11676] <= r_data[11675];
                
                r_data[11677] <= r_data[11676];
                
                r_data[11678] <= r_data[11677];
                
                r_data[11679] <= r_data[11678];
                
                r_data[11680] <= r_data[11679];
                
                r_data[11681] <= r_data[11680];
                
                r_data[11682] <= r_data[11681];
                
                r_data[11683] <= r_data[11682];
                
                r_data[11684] <= r_data[11683];
                
                r_data[11685] <= r_data[11684];
                
                r_data[11686] <= r_data[11685];
                
                r_data[11687] <= r_data[11686];
                
                r_data[11688] <= r_data[11687];
                
                r_data[11689] <= r_data[11688];
                
                r_data[11690] <= r_data[11689];
                
                r_data[11691] <= r_data[11690];
                
                r_data[11692] <= r_data[11691];
                
                r_data[11693] <= r_data[11692];
                
                r_data[11694] <= r_data[11693];
                
                r_data[11695] <= r_data[11694];
                
                r_data[11696] <= r_data[11695];
                
                r_data[11697] <= r_data[11696];
                
                r_data[11698] <= r_data[11697];
                
                r_data[11699] <= r_data[11698];
                
                r_data[11700] <= r_data[11699];
                
                r_data[11701] <= r_data[11700];
                
                r_data[11702] <= r_data[11701];
                
                r_data[11703] <= r_data[11702];
                
                r_data[11704] <= r_data[11703];
                
                r_data[11705] <= r_data[11704];
                
                r_data[11706] <= r_data[11705];
                
                r_data[11707] <= r_data[11706];
                
                r_data[11708] <= r_data[11707];
                
                r_data[11709] <= r_data[11708];
                
                r_data[11710] <= r_data[11709];
                
                r_data[11711] <= r_data[11710];
                
                r_data[11712] <= r_data[11711];
                
                r_data[11713] <= r_data[11712];
                
                r_data[11714] <= r_data[11713];
                
                r_data[11715] <= r_data[11714];
                
                r_data[11716] <= r_data[11715];
                
                r_data[11717] <= r_data[11716];
                
                r_data[11718] <= r_data[11717];
                
                r_data[11719] <= r_data[11718];
                
                r_data[11720] <= r_data[11719];
                
                r_data[11721] <= r_data[11720];
                
                r_data[11722] <= r_data[11721];
                
                r_data[11723] <= r_data[11722];
                
                r_data[11724] <= r_data[11723];
                
                r_data[11725] <= r_data[11724];
                
                r_data[11726] <= r_data[11725];
                
                r_data[11727] <= r_data[11726];
                
                r_data[11728] <= r_data[11727];
                
                r_data[11729] <= r_data[11728];
                
                r_data[11730] <= r_data[11729];
                
                r_data[11731] <= r_data[11730];
                
                r_data[11732] <= r_data[11731];
                
                r_data[11733] <= r_data[11732];
                
                r_data[11734] <= r_data[11733];
                
                r_data[11735] <= r_data[11734];
                
                r_data[11736] <= r_data[11735];
                
                r_data[11737] <= r_data[11736];
                
                r_data[11738] <= r_data[11737];
                
                r_data[11739] <= r_data[11738];
                
                r_data[11740] <= r_data[11739];
                
                r_data[11741] <= r_data[11740];
                
                r_data[11742] <= r_data[11741];
                
                r_data[11743] <= r_data[11742];
                
                r_data[11744] <= r_data[11743];
                
                r_data[11745] <= r_data[11744];
                
                r_data[11746] <= r_data[11745];
                
                r_data[11747] <= r_data[11746];
                
                r_data[11748] <= r_data[11747];
                
                r_data[11749] <= r_data[11748];
                
                r_data[11750] <= r_data[11749];
                
                r_data[11751] <= r_data[11750];
                
                r_data[11752] <= r_data[11751];
                
                r_data[11753] <= r_data[11752];
                
                r_data[11754] <= r_data[11753];
                
                r_data[11755] <= r_data[11754];
                
                r_data[11756] <= r_data[11755];
                
                r_data[11757] <= r_data[11756];
                
                r_data[11758] <= r_data[11757];
                
                r_data[11759] <= r_data[11758];
                
                r_data[11760] <= r_data[11759];
                
                r_data[11761] <= r_data[11760];
                
                r_data[11762] <= r_data[11761];
                
                r_data[11763] <= r_data[11762];
                
                r_data[11764] <= r_data[11763];
                
                r_data[11765] <= r_data[11764];
                
                r_data[11766] <= r_data[11765];
                
                r_data[11767] <= r_data[11766];
                
                r_data[11768] <= r_data[11767];
                
                r_data[11769] <= r_data[11768];
                
                r_data[11770] <= r_data[11769];
                
                r_data[11771] <= r_data[11770];
                
                r_data[11772] <= r_data[11771];
                
                r_data[11773] <= r_data[11772];
                
                r_data[11774] <= r_data[11773];
                
                r_data[11775] <= r_data[11774];
                
                r_data[11776] <= r_data[11775];
                
                r_data[11777] <= r_data[11776];
                
                r_data[11778] <= r_data[11777];
                
                r_data[11779] <= r_data[11778];
                
                r_data[11780] <= r_data[11779];
                
                r_data[11781] <= r_data[11780];
                
                r_data[11782] <= r_data[11781];
                
                r_data[11783] <= r_data[11782];
                
                r_data[11784] <= r_data[11783];
                
                r_data[11785] <= r_data[11784];
                
                r_data[11786] <= r_data[11785];
                
                r_data[11787] <= r_data[11786];
                
                r_data[11788] <= r_data[11787];
                
                r_data[11789] <= r_data[11788];
                
                r_data[11790] <= r_data[11789];
                
                r_data[11791] <= r_data[11790];
                
                r_data[11792] <= r_data[11791];
                
                r_data[11793] <= r_data[11792];
                
                r_data[11794] <= r_data[11793];
                
                r_data[11795] <= r_data[11794];
                
                r_data[11796] <= r_data[11795];
                
                r_data[11797] <= r_data[11796];
                
                r_data[11798] <= r_data[11797];
                
                r_data[11799] <= r_data[11798];
                
                r_data[11800] <= r_data[11799];
                
                r_data[11801] <= r_data[11800];
                
                r_data[11802] <= r_data[11801];
                
                r_data[11803] <= r_data[11802];
                
                r_data[11804] <= r_data[11803];
                
                r_data[11805] <= r_data[11804];
                
                r_data[11806] <= r_data[11805];
                
                r_data[11807] <= r_data[11806];
                
                r_data[11808] <= r_data[11807];
                
                r_data[11809] <= r_data[11808];
                
                r_data[11810] <= r_data[11809];
                
                r_data[11811] <= r_data[11810];
                
                r_data[11812] <= r_data[11811];
                
                r_data[11813] <= r_data[11812];
                
                r_data[11814] <= r_data[11813];
                
                r_data[11815] <= r_data[11814];
                
                r_data[11816] <= r_data[11815];
                
                r_data[11817] <= r_data[11816];
                
                r_data[11818] <= r_data[11817];
                
                r_data[11819] <= r_data[11818];
                
                r_data[11820] <= r_data[11819];
                
                r_data[11821] <= r_data[11820];
                
                r_data[11822] <= r_data[11821];
                
                r_data[11823] <= r_data[11822];
                
                r_data[11824] <= r_data[11823];
                
                r_data[11825] <= r_data[11824];
                
                r_data[11826] <= r_data[11825];
                
                r_data[11827] <= r_data[11826];
                
                r_data[11828] <= r_data[11827];
                
                r_data[11829] <= r_data[11828];
                
                r_data[11830] <= r_data[11829];
                
                r_data[11831] <= r_data[11830];
                
                r_data[11832] <= r_data[11831];
                
                r_data[11833] <= r_data[11832];
                
                r_data[11834] <= r_data[11833];
                
                r_data[11835] <= r_data[11834];
                
                r_data[11836] <= r_data[11835];
                
                r_data[11837] <= r_data[11836];
                
                r_data[11838] <= r_data[11837];
                
                r_data[11839] <= r_data[11838];
                
                r_data[11840] <= r_data[11839];
                
                r_data[11841] <= r_data[11840];
                
                r_data[11842] <= r_data[11841];
                
                r_data[11843] <= r_data[11842];
                
                r_data[11844] <= r_data[11843];
                
                r_data[11845] <= r_data[11844];
                
                r_data[11846] <= r_data[11845];
                
                r_data[11847] <= r_data[11846];
                
                r_data[11848] <= r_data[11847];
                
                r_data[11849] <= r_data[11848];
                
                r_data[11850] <= r_data[11849];
                
                r_data[11851] <= r_data[11850];
                
                r_data[11852] <= r_data[11851];
                
                r_data[11853] <= r_data[11852];
                
                r_data[11854] <= r_data[11853];
                
                r_data[11855] <= r_data[11854];
                
                r_data[11856] <= r_data[11855];
                
                r_data[11857] <= r_data[11856];
                
                r_data[11858] <= r_data[11857];
                
                r_data[11859] <= r_data[11858];
                
                r_data[11860] <= r_data[11859];
                
                r_data[11861] <= r_data[11860];
                
                r_data[11862] <= r_data[11861];
                
                r_data[11863] <= r_data[11862];
                
                r_data[11864] <= r_data[11863];
                
                r_data[11865] <= r_data[11864];
                
                r_data[11866] <= r_data[11865];
                
                r_data[11867] <= r_data[11866];
                
                r_data[11868] <= r_data[11867];
                
                r_data[11869] <= r_data[11868];
                
                r_data[11870] <= r_data[11869];
                
                r_data[11871] <= r_data[11870];
                
                r_data[11872] <= r_data[11871];
                
                r_data[11873] <= r_data[11872];
                
                r_data[11874] <= r_data[11873];
                
                r_data[11875] <= r_data[11874];
                
                r_data[11876] <= r_data[11875];
                
                r_data[11877] <= r_data[11876];
                
                r_data[11878] <= r_data[11877];
                
                r_data[11879] <= r_data[11878];
                
                r_data[11880] <= r_data[11879];
                
                r_data[11881] <= r_data[11880];
                
                r_data[11882] <= r_data[11881];
                
                r_data[11883] <= r_data[11882];
                
                r_data[11884] <= r_data[11883];
                
                r_data[11885] <= r_data[11884];
                
                r_data[11886] <= r_data[11885];
                
                r_data[11887] <= r_data[11886];
                
                r_data[11888] <= r_data[11887];
                
                r_data[11889] <= r_data[11888];
                
                r_data[11890] <= r_data[11889];
                
                r_data[11891] <= r_data[11890];
                
                r_data[11892] <= r_data[11891];
                
                r_data[11893] <= r_data[11892];
                
                r_data[11894] <= r_data[11893];
                
                r_data[11895] <= r_data[11894];
                
                r_data[11896] <= r_data[11895];
                
                r_data[11897] <= r_data[11896];
                
                r_data[11898] <= r_data[11897];
                
                r_data[11899] <= r_data[11898];
                
                r_data[11900] <= r_data[11899];
                
                r_data[11901] <= r_data[11900];
                
                r_data[11902] <= r_data[11901];
                
                r_data[11903] <= r_data[11902];
                
                r_data[11904] <= r_data[11903];
                
                r_data[11905] <= r_data[11904];
                
                r_data[11906] <= r_data[11905];
                
                r_data[11907] <= r_data[11906];
                
                r_data[11908] <= r_data[11907];
                
                r_data[11909] <= r_data[11908];
                
                r_data[11910] <= r_data[11909];
                
                r_data[11911] <= r_data[11910];
                
                r_data[11912] <= r_data[11911];
                
                r_data[11913] <= r_data[11912];
                
                r_data[11914] <= r_data[11913];
                
                r_data[11915] <= r_data[11914];
                
                r_data[11916] <= r_data[11915];
                
                r_data[11917] <= r_data[11916];
                
                r_data[11918] <= r_data[11917];
                
                r_data[11919] <= r_data[11918];
                
                r_data[11920] <= r_data[11919];
                
                r_data[11921] <= r_data[11920];
                
                r_data[11922] <= r_data[11921];
                
                r_data[11923] <= r_data[11922];
                
                r_data[11924] <= r_data[11923];
                
                r_data[11925] <= r_data[11924];
                
                r_data[11926] <= r_data[11925];
                
                r_data[11927] <= r_data[11926];
                
                r_data[11928] <= r_data[11927];
                
                r_data[11929] <= r_data[11928];
                
                r_data[11930] <= r_data[11929];
                
                r_data[11931] <= r_data[11930];
                
                r_data[11932] <= r_data[11931];
                
                r_data[11933] <= r_data[11932];
                
                r_data[11934] <= r_data[11933];
                
                r_data[11935] <= r_data[11934];
                
                r_data[11936] <= r_data[11935];
                
                r_data[11937] <= r_data[11936];
                
                r_data[11938] <= r_data[11937];
                
                r_data[11939] <= r_data[11938];
                
                r_data[11940] <= r_data[11939];
                
                r_data[11941] <= r_data[11940];
                
                r_data[11942] <= r_data[11941];
                
                r_data[11943] <= r_data[11942];
                
                r_data[11944] <= r_data[11943];
                
                r_data[11945] <= r_data[11944];
                
                r_data[11946] <= r_data[11945];
                
                r_data[11947] <= r_data[11946];
                
                r_data[11948] <= r_data[11947];
                
                r_data[11949] <= r_data[11948];
                
                r_data[11950] <= r_data[11949];
                
                r_data[11951] <= r_data[11950];
                
                r_data[11952] <= r_data[11951];
                
                r_data[11953] <= r_data[11952];
                
                r_data[11954] <= r_data[11953];
                
                r_data[11955] <= r_data[11954];
                
                r_data[11956] <= r_data[11955];
                
                r_data[11957] <= r_data[11956];
                
                r_data[11958] <= r_data[11957];
                
                r_data[11959] <= r_data[11958];
                
                r_data[11960] <= r_data[11959];
                
                r_data[11961] <= r_data[11960];
                
                r_data[11962] <= r_data[11961];
                
                r_data[11963] <= r_data[11962];
                
                r_data[11964] <= r_data[11963];
                
                r_data[11965] <= r_data[11964];
                
                r_data[11966] <= r_data[11965];
                
                r_data[11967] <= r_data[11966];
                
                r_data[11968] <= r_data[11967];
                
                r_data[11969] <= r_data[11968];
                
                r_data[11970] <= r_data[11969];
                
                r_data[11971] <= r_data[11970];
                
                r_data[11972] <= r_data[11971];
                
                r_data[11973] <= r_data[11972];
                
                r_data[11974] <= r_data[11973];
                
                r_data[11975] <= r_data[11974];
                
                r_data[11976] <= r_data[11975];
                
                r_data[11977] <= r_data[11976];
                
                r_data[11978] <= r_data[11977];
                
                r_data[11979] <= r_data[11978];
                
                r_data[11980] <= r_data[11979];
                
                r_data[11981] <= r_data[11980];
                
                r_data[11982] <= r_data[11981];
                
                r_data[11983] <= r_data[11982];
                
                r_data[11984] <= r_data[11983];
                
                r_data[11985] <= r_data[11984];
                
                r_data[11986] <= r_data[11985];
                
                r_data[11987] <= r_data[11986];
                
                r_data[11988] <= r_data[11987];
                
                r_data[11989] <= r_data[11988];
                
                r_data[11990] <= r_data[11989];
                
                r_data[11991] <= r_data[11990];
                
                r_data[11992] <= r_data[11991];
                
                r_data[11993] <= r_data[11992];
                
                r_data[11994] <= r_data[11993];
                
                r_data[11995] <= r_data[11994];
                
                r_data[11996] <= r_data[11995];
                
                r_data[11997] <= r_data[11996];
                
                r_data[11998] <= r_data[11997];
                
                r_data[11999] <= r_data[11998];
                
                r_data[12000] <= r_data[11999];
                
                r_data[12001] <= r_data[12000];
                
                r_data[12002] <= r_data[12001];
                
                r_data[12003] <= r_data[12002];
                
                r_data[12004] <= r_data[12003];
                
                r_data[12005] <= r_data[12004];
                
                r_data[12006] <= r_data[12005];
                
                r_data[12007] <= r_data[12006];
                
                r_data[12008] <= r_data[12007];
                
                r_data[12009] <= r_data[12008];
                
                r_data[12010] <= r_data[12009];
                
                r_data[12011] <= r_data[12010];
                
                r_data[12012] <= r_data[12011];
                
                r_data[12013] <= r_data[12012];
                
                r_data[12014] <= r_data[12013];
                
                r_data[12015] <= r_data[12014];
                
                r_data[12016] <= r_data[12015];
                
                r_data[12017] <= r_data[12016];
                
                r_data[12018] <= r_data[12017];
                
                r_data[12019] <= r_data[12018];
                
                r_data[12020] <= r_data[12019];
                
                r_data[12021] <= r_data[12020];
                
                r_data[12022] <= r_data[12021];
                
                r_data[12023] <= r_data[12022];
                
                r_data[12024] <= r_data[12023];
                
                r_data[12025] <= r_data[12024];
                
                r_data[12026] <= r_data[12025];
                
                r_data[12027] <= r_data[12026];
                
                r_data[12028] <= r_data[12027];
                
                r_data[12029] <= r_data[12028];
                
                r_data[12030] <= r_data[12029];
                
                r_data[12031] <= r_data[12030];
                
                r_data[12032] <= r_data[12031];
                
                r_data[12033] <= r_data[12032];
                
                r_data[12034] <= r_data[12033];
                
                r_data[12035] <= r_data[12034];
                
                r_data[12036] <= r_data[12035];
                
                r_data[12037] <= r_data[12036];
                
                r_data[12038] <= r_data[12037];
                
                r_data[12039] <= r_data[12038];
                
                r_data[12040] <= r_data[12039];
                
                r_data[12041] <= r_data[12040];
                
                r_data[12042] <= r_data[12041];
                
                r_data[12043] <= r_data[12042];
                
                r_data[12044] <= r_data[12043];
                
                r_data[12045] <= r_data[12044];
                
                r_data[12046] <= r_data[12045];
                
                r_data[12047] <= r_data[12046];
                
                r_data[12048] <= r_data[12047];
                
                r_data[12049] <= r_data[12048];
                
                r_data[12050] <= r_data[12049];
                
                r_data[12051] <= r_data[12050];
                
                r_data[12052] <= r_data[12051];
                
                r_data[12053] <= r_data[12052];
                
                r_data[12054] <= r_data[12053];
                
                r_data[12055] <= r_data[12054];
                
                r_data[12056] <= r_data[12055];
                
                r_data[12057] <= r_data[12056];
                
                r_data[12058] <= r_data[12057];
                
                r_data[12059] <= r_data[12058];
                
                r_data[12060] <= r_data[12059];
                
                r_data[12061] <= r_data[12060];
                
                r_data[12062] <= r_data[12061];
                
                r_data[12063] <= r_data[12062];
                
                r_data[12064] <= r_data[12063];
                
                r_data[12065] <= r_data[12064];
                
                r_data[12066] <= r_data[12065];
                
                r_data[12067] <= r_data[12066];
                
                r_data[12068] <= r_data[12067];
                
                r_data[12069] <= r_data[12068];
                
                r_data[12070] <= r_data[12069];
                
                r_data[12071] <= r_data[12070];
                
                r_data[12072] <= r_data[12071];
                
                r_data[12073] <= r_data[12072];
                
                r_data[12074] <= r_data[12073];
                
                r_data[12075] <= r_data[12074];
                
                r_data[12076] <= r_data[12075];
                
                r_data[12077] <= r_data[12076];
                
                r_data[12078] <= r_data[12077];
                
                r_data[12079] <= r_data[12078];
                
                r_data[12080] <= r_data[12079];
                
                r_data[12081] <= r_data[12080];
                
                r_data[12082] <= r_data[12081];
                
                r_data[12083] <= r_data[12082];
                
                r_data[12084] <= r_data[12083];
                
                r_data[12085] <= r_data[12084];
                
                r_data[12086] <= r_data[12085];
                
                r_data[12087] <= r_data[12086];
                
                r_data[12088] <= r_data[12087];
                
                r_data[12089] <= r_data[12088];
                
                r_data[12090] <= r_data[12089];
                
                r_data[12091] <= r_data[12090];
                
                r_data[12092] <= r_data[12091];
                
                r_data[12093] <= r_data[12092];
                
                r_data[12094] <= r_data[12093];
                
                r_data[12095] <= r_data[12094];
                
                r_data[12096] <= r_data[12095];
                
                r_data[12097] <= r_data[12096];
                
                r_data[12098] <= r_data[12097];
                
                r_data[12099] <= r_data[12098];
                
                r_data[12100] <= r_data[12099];
                
                r_data[12101] <= r_data[12100];
                
                r_data[12102] <= r_data[12101];
                
                r_data[12103] <= r_data[12102];
                
                r_data[12104] <= r_data[12103];
                
                r_data[12105] <= r_data[12104];
                
                r_data[12106] <= r_data[12105];
                
                r_data[12107] <= r_data[12106];
                
                r_data[12108] <= r_data[12107];
                
                r_data[12109] <= r_data[12108];
                
                r_data[12110] <= r_data[12109];
                
                r_data[12111] <= r_data[12110];
                
                r_data[12112] <= r_data[12111];
                
                r_data[12113] <= r_data[12112];
                
                r_data[12114] <= r_data[12113];
                
                r_data[12115] <= r_data[12114];
                
                r_data[12116] <= r_data[12115];
                
                r_data[12117] <= r_data[12116];
                
                r_data[12118] <= r_data[12117];
                
                r_data[12119] <= r_data[12118];
                
                r_data[12120] <= r_data[12119];
                
                r_data[12121] <= r_data[12120];
                
                r_data[12122] <= r_data[12121];
                
                r_data[12123] <= r_data[12122];
                
                r_data[12124] <= r_data[12123];
                
                r_data[12125] <= r_data[12124];
                
                r_data[12126] <= r_data[12125];
                
                r_data[12127] <= r_data[12126];
                
                r_data[12128] <= r_data[12127];
                
                r_data[12129] <= r_data[12128];
                
                r_data[12130] <= r_data[12129];
                
                r_data[12131] <= r_data[12130];
                
                r_data[12132] <= r_data[12131];
                
                r_data[12133] <= r_data[12132];
                
                r_data[12134] <= r_data[12133];
                
                r_data[12135] <= r_data[12134];
                
                r_data[12136] <= r_data[12135];
                
                r_data[12137] <= r_data[12136];
                
                r_data[12138] <= r_data[12137];
                
                r_data[12139] <= r_data[12138];
                
                r_data[12140] <= r_data[12139];
                
                r_data[12141] <= r_data[12140];
                
                r_data[12142] <= r_data[12141];
                
                r_data[12143] <= r_data[12142];
                
                r_data[12144] <= r_data[12143];
                
                r_data[12145] <= r_data[12144];
                
                r_data[12146] <= r_data[12145];
                
                r_data[12147] <= r_data[12146];
                
                r_data[12148] <= r_data[12147];
                
                r_data[12149] <= r_data[12148];
                
                r_data[12150] <= r_data[12149];
                
                r_data[12151] <= r_data[12150];
                
                r_data[12152] <= r_data[12151];
                
                r_data[12153] <= r_data[12152];
                
                r_data[12154] <= r_data[12153];
                
                r_data[12155] <= r_data[12154];
                
                r_data[12156] <= r_data[12155];
                
                r_data[12157] <= r_data[12156];
                
                r_data[12158] <= r_data[12157];
                
                r_data[12159] <= r_data[12158];
                
                r_data[12160] <= r_data[12159];
                
                r_data[12161] <= r_data[12160];
                
                r_data[12162] <= r_data[12161];
                
                r_data[12163] <= r_data[12162];
                
                r_data[12164] <= r_data[12163];
                
                r_data[12165] <= r_data[12164];
                
                r_data[12166] <= r_data[12165];
                
                r_data[12167] <= r_data[12166];
                
                r_data[12168] <= r_data[12167];
                
                r_data[12169] <= r_data[12168];
                
                r_data[12170] <= r_data[12169];
                
                r_data[12171] <= r_data[12170];
                
                r_data[12172] <= r_data[12171];
                
                r_data[12173] <= r_data[12172];
                
                r_data[12174] <= r_data[12173];
                
                r_data[12175] <= r_data[12174];
                
                r_data[12176] <= r_data[12175];
                
                r_data[12177] <= r_data[12176];
                
                r_data[12178] <= r_data[12177];
                
                r_data[12179] <= r_data[12178];
                
                r_data[12180] <= r_data[12179];
                
                r_data[12181] <= r_data[12180];
                
                r_data[12182] <= r_data[12181];
                
                r_data[12183] <= r_data[12182];
                
                r_data[12184] <= r_data[12183];
                
                r_data[12185] <= r_data[12184];
                
                r_data[12186] <= r_data[12185];
                
                r_data[12187] <= r_data[12186];
                
                r_data[12188] <= r_data[12187];
                
                r_data[12189] <= r_data[12188];
                
                r_data[12190] <= r_data[12189];
                
                r_data[12191] <= r_data[12190];
                
                r_data[12192] <= r_data[12191];
                
                r_data[12193] <= r_data[12192];
                
                r_data[12194] <= r_data[12193];
                
                r_data[12195] <= r_data[12194];
                
                r_data[12196] <= r_data[12195];
                
                r_data[12197] <= r_data[12196];
                
                r_data[12198] <= r_data[12197];
                
                r_data[12199] <= r_data[12198];
                
                r_data[12200] <= r_data[12199];
                
                r_data[12201] <= r_data[12200];
                
                r_data[12202] <= r_data[12201];
                
                r_data[12203] <= r_data[12202];
                
                r_data[12204] <= r_data[12203];
                
                r_data[12205] <= r_data[12204];
                
                r_data[12206] <= r_data[12205];
                
                r_data[12207] <= r_data[12206];
                
                r_data[12208] <= r_data[12207];
                
                r_data[12209] <= r_data[12208];
                
                r_data[12210] <= r_data[12209];
                
                r_data[12211] <= r_data[12210];
                
                r_data[12212] <= r_data[12211];
                
                r_data[12213] <= r_data[12212];
                
                r_data[12214] <= r_data[12213];
                
                r_data[12215] <= r_data[12214];
                
                r_data[12216] <= r_data[12215];
                
                r_data[12217] <= r_data[12216];
                
                r_data[12218] <= r_data[12217];
                
                r_data[12219] <= r_data[12218];
                
                r_data[12220] <= r_data[12219];
                
                r_data[12221] <= r_data[12220];
                
                r_data[12222] <= r_data[12221];
                
                r_data[12223] <= r_data[12222];
                
                r_data[12224] <= r_data[12223];
                
                r_data[12225] <= r_data[12224];
                
                r_data[12226] <= r_data[12225];
                
                r_data[12227] <= r_data[12226];
                
                r_data[12228] <= r_data[12227];
                
                r_data[12229] <= r_data[12228];
                
                r_data[12230] <= r_data[12229];
                
                r_data[12231] <= r_data[12230];
                
                r_data[12232] <= r_data[12231];
                
                r_data[12233] <= r_data[12232];
                
                r_data[12234] <= r_data[12233];
                
                r_data[12235] <= r_data[12234];
                
                r_data[12236] <= r_data[12235];
                
                r_data[12237] <= r_data[12236];
                
                r_data[12238] <= r_data[12237];
                
                r_data[12239] <= r_data[12238];
                
                r_data[12240] <= r_data[12239];
                
                r_data[12241] <= r_data[12240];
                
                r_data[12242] <= r_data[12241];
                
                r_data[12243] <= r_data[12242];
                
                r_data[12244] <= r_data[12243];
                
                r_data[12245] <= r_data[12244];
                
                r_data[12246] <= r_data[12245];
                
                r_data[12247] <= r_data[12246];
                
                r_data[12248] <= r_data[12247];
                
                r_data[12249] <= r_data[12248];
                
                r_data[12250] <= r_data[12249];
                
                r_data[12251] <= r_data[12250];
                
                r_data[12252] <= r_data[12251];
                
                r_data[12253] <= r_data[12252];
                
                r_data[12254] <= r_data[12253];
                
                r_data[12255] <= r_data[12254];
                
                r_data[12256] <= r_data[12255];
                
                r_data[12257] <= r_data[12256];
                
                r_data[12258] <= r_data[12257];
                
                r_data[12259] <= r_data[12258];
                
                r_data[12260] <= r_data[12259];
                
                r_data[12261] <= r_data[12260];
                
                r_data[12262] <= r_data[12261];
                
                r_data[12263] <= r_data[12262];
                
                r_data[12264] <= r_data[12263];
                
                r_data[12265] <= r_data[12264];
                
                r_data[12266] <= r_data[12265];
                
                r_data[12267] <= r_data[12266];
                
                r_data[12268] <= r_data[12267];
                
                r_data[12269] <= r_data[12268];
                
                r_data[12270] <= r_data[12269];
                
                r_data[12271] <= r_data[12270];
                
                r_data[12272] <= r_data[12271];
                
                r_data[12273] <= r_data[12272];
                
                r_data[12274] <= r_data[12273];
                
                r_data[12275] <= r_data[12274];
                
                r_data[12276] <= r_data[12275];
                
                r_data[12277] <= r_data[12276];
                
                r_data[12278] <= r_data[12277];
                
                r_data[12279] <= r_data[12278];
                
                r_data[12280] <= r_data[12279];
                
                r_data[12281] <= r_data[12280];
                
                r_data[12282] <= r_data[12281];
                
                r_data[12283] <= r_data[12282];
                
                r_data[12284] <= r_data[12283];
                
                r_data[12285] <= r_data[12284];
                
                r_data[12286] <= r_data[12285];
                
                r_data[12287] <= r_data[12286];
                
                r_data[12288] <= r_data[12287];
                
                r_data[12289] <= r_data[12288];
                
                r_data[12290] <= r_data[12289];
                
                r_data[12291] <= r_data[12290];
                
                r_data[12292] <= r_data[12291];
                
                r_data[12293] <= r_data[12292];
                
                r_data[12294] <= r_data[12293];
                
                r_data[12295] <= r_data[12294];
                
                r_data[12296] <= r_data[12295];
                
                r_data[12297] <= r_data[12296];
                
                r_data[12298] <= r_data[12297];
                
                r_data[12299] <= r_data[12298];
                
                r_data[12300] <= r_data[12299];
                
                r_data[12301] <= r_data[12300];
                
                r_data[12302] <= r_data[12301];
                
                r_data[12303] <= r_data[12302];
                
                r_data[12304] <= r_data[12303];
                
                r_data[12305] <= r_data[12304];
                
                r_data[12306] <= r_data[12305];
                
                r_data[12307] <= r_data[12306];
                
                r_data[12308] <= r_data[12307];
                
                r_data[12309] <= r_data[12308];
                
                r_data[12310] <= r_data[12309];
                
                r_data[12311] <= r_data[12310];
                
                r_data[12312] <= r_data[12311];
                
                r_data[12313] <= r_data[12312];
                
                r_data[12314] <= r_data[12313];
                
                r_data[12315] <= r_data[12314];
                
                r_data[12316] <= r_data[12315];
                
                r_data[12317] <= r_data[12316];
                
                r_data[12318] <= r_data[12317];
                
                r_data[12319] <= r_data[12318];
                
                r_data[12320] <= r_data[12319];
                
                r_data[12321] <= r_data[12320];
                
                r_data[12322] <= r_data[12321];
                
                r_data[12323] <= r_data[12322];
                
                r_data[12324] <= r_data[12323];
                
                r_data[12325] <= r_data[12324];
                
                r_data[12326] <= r_data[12325];
                
                r_data[12327] <= r_data[12326];
                
                r_data[12328] <= r_data[12327];
                
                r_data[12329] <= r_data[12328];
                
                r_data[12330] <= r_data[12329];
                
                r_data[12331] <= r_data[12330];
                
                r_data[12332] <= r_data[12331];
                
                r_data[12333] <= r_data[12332];
                
                r_data[12334] <= r_data[12333];
                
                r_data[12335] <= r_data[12334];
                
                r_data[12336] <= r_data[12335];
                
                r_data[12337] <= r_data[12336];
                
                r_data[12338] <= r_data[12337];
                
                r_data[12339] <= r_data[12338];
                
                r_data[12340] <= r_data[12339];
                
                r_data[12341] <= r_data[12340];
                
                r_data[12342] <= r_data[12341];
                
                r_data[12343] <= r_data[12342];
                
                r_data[12344] <= r_data[12343];
                
                r_data[12345] <= r_data[12344];
                
                r_data[12346] <= r_data[12345];
                
                r_data[12347] <= r_data[12346];
                
                r_data[12348] <= r_data[12347];
                
                r_data[12349] <= r_data[12348];
                
                r_data[12350] <= r_data[12349];
                
                r_data[12351] <= r_data[12350];
                
                r_data[12352] <= r_data[12351];
                
                r_data[12353] <= r_data[12352];
                
                r_data[12354] <= r_data[12353];
                
                r_data[12355] <= r_data[12354];
                
                r_data[12356] <= r_data[12355];
                
                r_data[12357] <= r_data[12356];
                
                r_data[12358] <= r_data[12357];
                
                r_data[12359] <= r_data[12358];
                
                r_data[12360] <= r_data[12359];
                
                r_data[12361] <= r_data[12360];
                
                r_data[12362] <= r_data[12361];
                
                r_data[12363] <= r_data[12362];
                
                r_data[12364] <= r_data[12363];
                
                r_data[12365] <= r_data[12364];
                
                r_data[12366] <= r_data[12365];
                
                r_data[12367] <= r_data[12366];
                
                r_data[12368] <= r_data[12367];
                
                r_data[12369] <= r_data[12368];
                
                r_data[12370] <= r_data[12369];
                
                r_data[12371] <= r_data[12370];
                
                r_data[12372] <= r_data[12371];
                
                r_data[12373] <= r_data[12372];
                
                r_data[12374] <= r_data[12373];
                
                r_data[12375] <= r_data[12374];
                
                r_data[12376] <= r_data[12375];
                
                r_data[12377] <= r_data[12376];
                
                r_data[12378] <= r_data[12377];
                
                r_data[12379] <= r_data[12378];
                
                r_data[12380] <= r_data[12379];
                
                r_data[12381] <= r_data[12380];
                
                r_data[12382] <= r_data[12381];
                
                r_data[12383] <= r_data[12382];
                
                r_data[12384] <= r_data[12383];
                
                r_data[12385] <= r_data[12384];
                
                r_data[12386] <= r_data[12385];
                
                r_data[12387] <= r_data[12386];
                
                r_data[12388] <= r_data[12387];
                
                r_data[12389] <= r_data[12388];
                
                r_data[12390] <= r_data[12389];
                
                r_data[12391] <= r_data[12390];
                
                r_data[12392] <= r_data[12391];
                
                r_data[12393] <= r_data[12392];
                
                r_data[12394] <= r_data[12393];
                
                r_data[12395] <= r_data[12394];
                
                r_data[12396] <= r_data[12395];
                
                r_data[12397] <= r_data[12396];
                
                r_data[12398] <= r_data[12397];
                
                r_data[12399] <= r_data[12398];
                
                r_data[12400] <= r_data[12399];
                
                r_data[12401] <= r_data[12400];
                
                r_data[12402] <= r_data[12401];
                
                r_data[12403] <= r_data[12402];
                
                r_data[12404] <= r_data[12403];
                
                r_data[12405] <= r_data[12404];
                
                r_data[12406] <= r_data[12405];
                
                r_data[12407] <= r_data[12406];
                
                r_data[12408] <= r_data[12407];
                
                r_data[12409] <= r_data[12408];
                
                r_data[12410] <= r_data[12409];
                
                r_data[12411] <= r_data[12410];
                
                r_data[12412] <= r_data[12411];
                
                r_data[12413] <= r_data[12412];
                
                r_data[12414] <= r_data[12413];
                
                r_data[12415] <= r_data[12414];
                
                r_data[12416] <= r_data[12415];
                
                r_data[12417] <= r_data[12416];
                
                r_data[12418] <= r_data[12417];
                
                r_data[12419] <= r_data[12418];
                
                r_data[12420] <= r_data[12419];
                
                r_data[12421] <= r_data[12420];
                
                r_data[12422] <= r_data[12421];
                
                r_data[12423] <= r_data[12422];
                
                r_data[12424] <= r_data[12423];
                
                r_data[12425] <= r_data[12424];
                
                r_data[12426] <= r_data[12425];
                
                r_data[12427] <= r_data[12426];
                
                r_data[12428] <= r_data[12427];
                
                r_data[12429] <= r_data[12428];
                
                r_data[12430] <= r_data[12429];
                
                r_data[12431] <= r_data[12430];
                
                r_data[12432] <= r_data[12431];
                
                r_data[12433] <= r_data[12432];
                
                r_data[12434] <= r_data[12433];
                
                r_data[12435] <= r_data[12434];
                
                r_data[12436] <= r_data[12435];
                
                r_data[12437] <= r_data[12436];
                
                r_data[12438] <= r_data[12437];
                
                r_data[12439] <= r_data[12438];
                
                r_data[12440] <= r_data[12439];
                
                r_data[12441] <= r_data[12440];
                
                r_data[12442] <= r_data[12441];
                
                r_data[12443] <= r_data[12442];
                
                r_data[12444] <= r_data[12443];
                
                r_data[12445] <= r_data[12444];
                
                r_data[12446] <= r_data[12445];
                
                r_data[12447] <= r_data[12446];
                
                r_data[12448] <= r_data[12447];
                
                r_data[12449] <= r_data[12448];
                
                r_data[12450] <= r_data[12449];
                
                r_data[12451] <= r_data[12450];
                
                r_data[12452] <= r_data[12451];
                
                r_data[12453] <= r_data[12452];
                
                r_data[12454] <= r_data[12453];
                
                r_data[12455] <= r_data[12454];
                
                r_data[12456] <= r_data[12455];
                
                r_data[12457] <= r_data[12456];
                
                r_data[12458] <= r_data[12457];
                
                r_data[12459] <= r_data[12458];
                
                r_data[12460] <= r_data[12459];
                
                r_data[12461] <= r_data[12460];
                
                r_data[12462] <= r_data[12461];
                
                r_data[12463] <= r_data[12462];
                
                r_data[12464] <= r_data[12463];
                
                r_data[12465] <= r_data[12464];
                
                r_data[12466] <= r_data[12465];
                
                r_data[12467] <= r_data[12466];
                
                r_data[12468] <= r_data[12467];
                
                r_data[12469] <= r_data[12468];
                
                r_data[12470] <= r_data[12469];
                
                r_data[12471] <= r_data[12470];
                
                r_data[12472] <= r_data[12471];
                
                r_data[12473] <= r_data[12472];
                
                r_data[12474] <= r_data[12473];
                
                r_data[12475] <= r_data[12474];
                
                r_data[12476] <= r_data[12475];
                
                r_data[12477] <= r_data[12476];
                
                r_data[12478] <= r_data[12477];
                
                r_data[12479] <= r_data[12478];
                
                r_data[12480] <= r_data[12479];
                
                r_data[12481] <= r_data[12480];
                
                r_data[12482] <= r_data[12481];
                
                r_data[12483] <= r_data[12482];
                
                r_data[12484] <= r_data[12483];
                
                r_data[12485] <= r_data[12484];
                
                r_data[12486] <= r_data[12485];
                
                r_data[12487] <= r_data[12486];
                
                r_data[12488] <= r_data[12487];
                
                r_data[12489] <= r_data[12488];
                
                r_data[12490] <= r_data[12489];
                
                r_data[12491] <= r_data[12490];
                
                r_data[12492] <= r_data[12491];
                
                r_data[12493] <= r_data[12492];
                
                r_data[12494] <= r_data[12493];
                
                r_data[12495] <= r_data[12494];
                
                r_data[12496] <= r_data[12495];
                
                r_data[12497] <= r_data[12496];
                
                r_data[12498] <= r_data[12497];
                
                r_data[12499] <= r_data[12498];
                
                r_data[12500] <= r_data[12499];
                
                r_data[12501] <= r_data[12500];
                
                r_data[12502] <= r_data[12501];
                
                r_data[12503] <= r_data[12502];
                
                r_data[12504] <= r_data[12503];
                
                r_data[12505] <= r_data[12504];
                
                r_data[12506] <= r_data[12505];
                
                r_data[12507] <= r_data[12506];
                
                r_data[12508] <= r_data[12507];
                
                r_data[12509] <= r_data[12508];
                
                r_data[12510] <= r_data[12509];
                
                r_data[12511] <= r_data[12510];
                
                r_data[12512] <= r_data[12511];
                
                r_data[12513] <= r_data[12512];
                
                r_data[12514] <= r_data[12513];
                
                r_data[12515] <= r_data[12514];
                
                r_data[12516] <= r_data[12515];
                
                r_data[12517] <= r_data[12516];
                
                r_data[12518] <= r_data[12517];
                
                r_data[12519] <= r_data[12518];
                
                r_data[12520] <= r_data[12519];
                
                r_data[12521] <= r_data[12520];
                
                r_data[12522] <= r_data[12521];
                
                r_data[12523] <= r_data[12522];
                
                r_data[12524] <= r_data[12523];
                
                r_data[12525] <= r_data[12524];
                
                r_data[12526] <= r_data[12525];
                
                r_data[12527] <= r_data[12526];
                
                r_data[12528] <= r_data[12527];
                
                r_data[12529] <= r_data[12528];
                
                r_data[12530] <= r_data[12529];
                
                r_data[12531] <= r_data[12530];
                
                r_data[12532] <= r_data[12531];
                
                r_data[12533] <= r_data[12532];
                
                r_data[12534] <= r_data[12533];
                
                r_data[12535] <= r_data[12534];
                
                r_data[12536] <= r_data[12535];
                
                r_data[12537] <= r_data[12536];
                
                r_data[12538] <= r_data[12537];
                
                r_data[12539] <= r_data[12538];
                
                r_data[12540] <= r_data[12539];
                
                r_data[12541] <= r_data[12540];
                
                r_data[12542] <= r_data[12541];
                
                r_data[12543] <= r_data[12542];
                
                r_data[12544] <= r_data[12543];
                
                r_data[12545] <= r_data[12544];
                
                r_data[12546] <= r_data[12545];
                
                r_data[12547] <= r_data[12546];
                
                r_data[12548] <= r_data[12547];
                
                r_data[12549] <= r_data[12548];
                
                r_data[12550] <= r_data[12549];
                
                r_data[12551] <= r_data[12550];
                
                r_data[12552] <= r_data[12551];
                
                r_data[12553] <= r_data[12552];
                
                r_data[12554] <= r_data[12553];
                
                r_data[12555] <= r_data[12554];
                
                r_data[12556] <= r_data[12555];
                
                r_data[12557] <= r_data[12556];
                
                r_data[12558] <= r_data[12557];
                
                r_data[12559] <= r_data[12558];
                
                r_data[12560] <= r_data[12559];
                
                r_data[12561] <= r_data[12560];
                
                r_data[12562] <= r_data[12561];
                
                r_data[12563] <= r_data[12562];
                
                r_data[12564] <= r_data[12563];
                
                r_data[12565] <= r_data[12564];
                
                r_data[12566] <= r_data[12565];
                
                r_data[12567] <= r_data[12566];
                
                r_data[12568] <= r_data[12567];
                
                r_data[12569] <= r_data[12568];
                
                r_data[12570] <= r_data[12569];
                
                r_data[12571] <= r_data[12570];
                
                r_data[12572] <= r_data[12571];
                
                r_data[12573] <= r_data[12572];
                
                r_data[12574] <= r_data[12573];
                
                r_data[12575] <= r_data[12574];
                
                r_data[12576] <= r_data[12575];
                
                r_data[12577] <= r_data[12576];
                
                r_data[12578] <= r_data[12577];
                
                r_data[12579] <= r_data[12578];
                
                r_data[12580] <= r_data[12579];
                
                r_data[12581] <= r_data[12580];
                
                r_data[12582] <= r_data[12581];
                
                r_data[12583] <= r_data[12582];
                
                r_data[12584] <= r_data[12583];
                
                r_data[12585] <= r_data[12584];
                
                r_data[12586] <= r_data[12585];
                
                r_data[12587] <= r_data[12586];
                
                r_data[12588] <= r_data[12587];
                
                r_data[12589] <= r_data[12588];
                
                r_data[12590] <= r_data[12589];
                
                r_data[12591] <= r_data[12590];
                
                r_data[12592] <= r_data[12591];
                
                r_data[12593] <= r_data[12592];
                
                r_data[12594] <= r_data[12593];
                
                r_data[12595] <= r_data[12594];
                
                r_data[12596] <= r_data[12595];
                
                r_data[12597] <= r_data[12596];
                
                r_data[12598] <= r_data[12597];
                
                r_data[12599] <= r_data[12598];
                
                r_data[12600] <= r_data[12599];
                
                r_data[12601] <= r_data[12600];
                
                r_data[12602] <= r_data[12601];
                
                r_data[12603] <= r_data[12602];
                
                r_data[12604] <= r_data[12603];
                
                r_data[12605] <= r_data[12604];
                
                r_data[12606] <= r_data[12605];
                
                r_data[12607] <= r_data[12606];
                
                r_data[12608] <= r_data[12607];
                
                r_data[12609] <= r_data[12608];
                
                r_data[12610] <= r_data[12609];
                
                r_data[12611] <= r_data[12610];
                
                r_data[12612] <= r_data[12611];
                
                r_data[12613] <= r_data[12612];
                
                r_data[12614] <= r_data[12613];
                
                r_data[12615] <= r_data[12614];
                
                r_data[12616] <= r_data[12615];
                
                r_data[12617] <= r_data[12616];
                
                r_data[12618] <= r_data[12617];
                
                r_data[12619] <= r_data[12618];
                
                r_data[12620] <= r_data[12619];
                
                r_data[12621] <= r_data[12620];
                
                r_data[12622] <= r_data[12621];
                
                r_data[12623] <= r_data[12622];
                
                r_data[12624] <= r_data[12623];
                
                r_data[12625] <= r_data[12624];
                
                r_data[12626] <= r_data[12625];
                
                r_data[12627] <= r_data[12626];
                
                r_data[12628] <= r_data[12627];
                
                r_data[12629] <= r_data[12628];
                
                r_data[12630] <= r_data[12629];
                
                r_data[12631] <= r_data[12630];
                
                r_data[12632] <= r_data[12631];
                
                r_data[12633] <= r_data[12632];
                
                r_data[12634] <= r_data[12633];
                
                r_data[12635] <= r_data[12634];
                
                r_data[12636] <= r_data[12635];
                
                r_data[12637] <= r_data[12636];
                
                r_data[12638] <= r_data[12637];
                
                r_data[12639] <= r_data[12638];
                
                r_data[12640] <= r_data[12639];
                
                r_data[12641] <= r_data[12640];
                
                r_data[12642] <= r_data[12641];
                
                r_data[12643] <= r_data[12642];
                
                r_data[12644] <= r_data[12643];
                
                r_data[12645] <= r_data[12644];
                
                r_data[12646] <= r_data[12645];
                
                r_data[12647] <= r_data[12646];
                
                r_data[12648] <= r_data[12647];
                
                r_data[12649] <= r_data[12648];
                
                r_data[12650] <= r_data[12649];
                
                r_data[12651] <= r_data[12650];
                
                r_data[12652] <= r_data[12651];
                
                r_data[12653] <= r_data[12652];
                
                r_data[12654] <= r_data[12653];
                
                r_data[12655] <= r_data[12654];
                
                r_data[12656] <= r_data[12655];
                
                r_data[12657] <= r_data[12656];
                
                r_data[12658] <= r_data[12657];
                
                r_data[12659] <= r_data[12658];
                
                r_data[12660] <= r_data[12659];
                
                r_data[12661] <= r_data[12660];
                
                r_data[12662] <= r_data[12661];
                
                r_data[12663] <= r_data[12662];
                
                r_data[12664] <= r_data[12663];
                
                r_data[12665] <= r_data[12664];
                
                r_data[12666] <= r_data[12665];
                
                r_data[12667] <= r_data[12666];
                
                r_data[12668] <= r_data[12667];
                
                r_data[12669] <= r_data[12668];
                
                r_data[12670] <= r_data[12669];
                
                r_data[12671] <= r_data[12670];
                
                r_data[12672] <= r_data[12671];
                
                r_data[12673] <= r_data[12672];
                
                r_data[12674] <= r_data[12673];
                
                r_data[12675] <= r_data[12674];
                
                r_data[12676] <= r_data[12675];
                
                r_data[12677] <= r_data[12676];
                
                r_data[12678] <= r_data[12677];
                
                r_data[12679] <= r_data[12678];
                
                r_data[12680] <= r_data[12679];
                
                r_data[12681] <= r_data[12680];
                
                r_data[12682] <= r_data[12681];
                
                r_data[12683] <= r_data[12682];
                
                r_data[12684] <= r_data[12683];
                
                r_data[12685] <= r_data[12684];
                
                r_data[12686] <= r_data[12685];
                
                r_data[12687] <= r_data[12686];
                
                r_data[12688] <= r_data[12687];
                
                r_data[12689] <= r_data[12688];
                
                r_data[12690] <= r_data[12689];
                
                r_data[12691] <= r_data[12690];
                
                r_data[12692] <= r_data[12691];
                
                r_data[12693] <= r_data[12692];
                
                r_data[12694] <= r_data[12693];
                
                r_data[12695] <= r_data[12694];
                
                r_data[12696] <= r_data[12695];
                
                r_data[12697] <= r_data[12696];
                
                r_data[12698] <= r_data[12697];
                
                r_data[12699] <= r_data[12698];
                
                r_data[12700] <= r_data[12699];
                
                r_data[12701] <= r_data[12700];
                
                r_data[12702] <= r_data[12701];
                
                r_data[12703] <= r_data[12702];
                
                r_data[12704] <= r_data[12703];
                
                r_data[12705] <= r_data[12704];
                
                r_data[12706] <= r_data[12705];
                
                r_data[12707] <= r_data[12706];
                
                r_data[12708] <= r_data[12707];
                
                r_data[12709] <= r_data[12708];
                
                r_data[12710] <= r_data[12709];
                
                r_data[12711] <= r_data[12710];
                
                r_data[12712] <= r_data[12711];
                
                r_data[12713] <= r_data[12712];
                
                r_data[12714] <= r_data[12713];
                
                r_data[12715] <= r_data[12714];
                
                r_data[12716] <= r_data[12715];
                
                r_data[12717] <= r_data[12716];
                
                r_data[12718] <= r_data[12717];
                
                r_data[12719] <= r_data[12718];
                
                r_data[12720] <= r_data[12719];
                
                r_data[12721] <= r_data[12720];
                
                r_data[12722] <= r_data[12721];
                
                r_data[12723] <= r_data[12722];
                
                r_data[12724] <= r_data[12723];
                
                r_data[12725] <= r_data[12724];
                
                r_data[12726] <= r_data[12725];
                
                r_data[12727] <= r_data[12726];
                
                r_data[12728] <= r_data[12727];
                
                r_data[12729] <= r_data[12728];
                
                r_data[12730] <= r_data[12729];
                
                r_data[12731] <= r_data[12730];
                
                r_data[12732] <= r_data[12731];
                
                r_data[12733] <= r_data[12732];
                
                r_data[12734] <= r_data[12733];
                
                r_data[12735] <= r_data[12734];
                
                r_data[12736] <= r_data[12735];
                
                r_data[12737] <= r_data[12736];
                
                r_data[12738] <= r_data[12737];
                
                r_data[12739] <= r_data[12738];
                
                r_data[12740] <= r_data[12739];
                
                r_data[12741] <= r_data[12740];
                
                r_data[12742] <= r_data[12741];
                
                r_data[12743] <= r_data[12742];
                
                r_data[12744] <= r_data[12743];
                
                r_data[12745] <= r_data[12744];
                
                r_data[12746] <= r_data[12745];
                
                r_data[12747] <= r_data[12746];
                
                r_data[12748] <= r_data[12747];
                
                r_data[12749] <= r_data[12748];
                
                r_data[12750] <= r_data[12749];
                
                r_data[12751] <= r_data[12750];
                
                r_data[12752] <= r_data[12751];
                
                r_data[12753] <= r_data[12752];
                
                r_data[12754] <= r_data[12753];
                
                r_data[12755] <= r_data[12754];
                
                r_data[12756] <= r_data[12755];
                
                r_data[12757] <= r_data[12756];
                
                r_data[12758] <= r_data[12757];
                
                r_data[12759] <= r_data[12758];
                
                r_data[12760] <= r_data[12759];
                
                r_data[12761] <= r_data[12760];
                
                r_data[12762] <= r_data[12761];
                
                r_data[12763] <= r_data[12762];
                
                r_data[12764] <= r_data[12763];
                
                r_data[12765] <= r_data[12764];
                
                r_data[12766] <= r_data[12765];
                
                r_data[12767] <= r_data[12766];
                
                r_data[12768] <= r_data[12767];
                
                r_data[12769] <= r_data[12768];
                
                r_data[12770] <= r_data[12769];
                
                r_data[12771] <= r_data[12770];
                
                r_data[12772] <= r_data[12771];
                
                r_data[12773] <= r_data[12772];
                
                r_data[12774] <= r_data[12773];
                
                r_data[12775] <= r_data[12774];
                
                r_data[12776] <= r_data[12775];
                
                r_data[12777] <= r_data[12776];
                
                r_data[12778] <= r_data[12777];
                
                r_data[12779] <= r_data[12778];
                
                r_data[12780] <= r_data[12779];
                
                r_data[12781] <= r_data[12780];
                
                r_data[12782] <= r_data[12781];
                
                r_data[12783] <= r_data[12782];
                
                r_data[12784] <= r_data[12783];
                
                r_data[12785] <= r_data[12784];
                
                r_data[12786] <= r_data[12785];
                
                r_data[12787] <= r_data[12786];
                
                r_data[12788] <= r_data[12787];
                
                r_data[12789] <= r_data[12788];
                
                r_data[12790] <= r_data[12789];
                
                r_data[12791] <= r_data[12790];
                
                r_data[12792] <= r_data[12791];
                
                r_data[12793] <= r_data[12792];
                
                r_data[12794] <= r_data[12793];
                
                r_data[12795] <= r_data[12794];
                
                r_data[12796] <= r_data[12795];
                
                r_data[12797] <= r_data[12796];
                
                r_data[12798] <= r_data[12797];
                
                r_data[12799] <= r_data[12798];
                
                r_data[12800] <= r_data[12799];
                
                r_data[12801] <= r_data[12800];
                
                r_data[12802] <= r_data[12801];
                
                r_data[12803] <= r_data[12802];
                
                r_data[12804] <= r_data[12803];
                
                r_data[12805] <= r_data[12804];
                
                r_data[12806] <= r_data[12805];
                
                r_data[12807] <= r_data[12806];
                
                r_data[12808] <= r_data[12807];
                
                r_data[12809] <= r_data[12808];
                
                r_data[12810] <= r_data[12809];
                
                r_data[12811] <= r_data[12810];
                
                r_data[12812] <= r_data[12811];
                
                r_data[12813] <= r_data[12812];
                
                r_data[12814] <= r_data[12813];
                
                r_data[12815] <= r_data[12814];
                
                r_data[12816] <= r_data[12815];
                
                r_data[12817] <= r_data[12816];
                
                r_data[12818] <= r_data[12817];
                
                r_data[12819] <= r_data[12818];
                
                r_data[12820] <= r_data[12819];
                
                r_data[12821] <= r_data[12820];
                
                r_data[12822] <= r_data[12821];
                
                r_data[12823] <= r_data[12822];
                
                r_data[12824] <= r_data[12823];
                
                r_data[12825] <= r_data[12824];
                
                r_data[12826] <= r_data[12825];
                
                r_data[12827] <= r_data[12826];
                
                r_data[12828] <= r_data[12827];
                
                r_data[12829] <= r_data[12828];
                
                r_data[12830] <= r_data[12829];
                
                r_data[12831] <= r_data[12830];
                
                r_data[12832] <= r_data[12831];
                
                r_data[12833] <= r_data[12832];
                
                r_data[12834] <= r_data[12833];
                
                r_data[12835] <= r_data[12834];
                
                r_data[12836] <= r_data[12835];
                
                r_data[12837] <= r_data[12836];
                
                r_data[12838] <= r_data[12837];
                
                r_data[12839] <= r_data[12838];
                
                r_data[12840] <= r_data[12839];
                
                r_data[12841] <= r_data[12840];
                
                r_data[12842] <= r_data[12841];
                
                r_data[12843] <= r_data[12842];
                
                r_data[12844] <= r_data[12843];
                
                r_data[12845] <= r_data[12844];
                
                r_data[12846] <= r_data[12845];
                
                r_data[12847] <= r_data[12846];
                
                r_data[12848] <= r_data[12847];
                
                r_data[12849] <= r_data[12848];
                
                r_data[12850] <= r_data[12849];
                
                r_data[12851] <= r_data[12850];
                
                r_data[12852] <= r_data[12851];
                
                r_data[12853] <= r_data[12852];
                
                r_data[12854] <= r_data[12853];
                
                r_data[12855] <= r_data[12854];
                
                r_data[12856] <= r_data[12855];
                
                r_data[12857] <= r_data[12856];
                
                r_data[12858] <= r_data[12857];
                
                r_data[12859] <= r_data[12858];
                
                r_data[12860] <= r_data[12859];
                
                r_data[12861] <= r_data[12860];
                
                r_data[12862] <= r_data[12861];
                
                r_data[12863] <= r_data[12862];
                
                r_data[12864] <= r_data[12863];
                
                r_data[12865] <= r_data[12864];
                
                r_data[12866] <= r_data[12865];
                
                r_data[12867] <= r_data[12866];
                
                r_data[12868] <= r_data[12867];
                
                r_data[12869] <= r_data[12868];
                
                r_data[12870] <= r_data[12869];
                
                r_data[12871] <= r_data[12870];
                
                r_data[12872] <= r_data[12871];
                
                r_data[12873] <= r_data[12872];
                
                r_data[12874] <= r_data[12873];
                
                r_data[12875] <= r_data[12874];
                
                r_data[12876] <= r_data[12875];
                
                r_data[12877] <= r_data[12876];
                
                r_data[12878] <= r_data[12877];
                
                r_data[12879] <= r_data[12878];
                
                r_data[12880] <= r_data[12879];
                
                r_data[12881] <= r_data[12880];
                
                r_data[12882] <= r_data[12881];
                
                r_data[12883] <= r_data[12882];
                
                r_data[12884] <= r_data[12883];
                
                r_data[12885] <= r_data[12884];
                
                r_data[12886] <= r_data[12885];
                
                r_data[12887] <= r_data[12886];
                
                r_data[12888] <= r_data[12887];
                
                r_data[12889] <= r_data[12888];
                
                r_data[12890] <= r_data[12889];
                
                r_data[12891] <= r_data[12890];
                
                r_data[12892] <= r_data[12891];
                
                r_data[12893] <= r_data[12892];
                
                r_data[12894] <= r_data[12893];
                
                r_data[12895] <= r_data[12894];
                
                r_data[12896] <= r_data[12895];
                
                r_data[12897] <= r_data[12896];
                
                r_data[12898] <= r_data[12897];
                
                r_data[12899] <= r_data[12898];
                
                r_data[12900] <= r_data[12899];
                
                r_data[12901] <= r_data[12900];
                
                r_data[12902] <= r_data[12901];
                
                r_data[12903] <= r_data[12902];
                
                r_data[12904] <= r_data[12903];
                
                r_data[12905] <= r_data[12904];
                
                r_data[12906] <= r_data[12905];
                
                r_data[12907] <= r_data[12906];
                
                r_data[12908] <= r_data[12907];
                
                r_data[12909] <= r_data[12908];
                
                r_data[12910] <= r_data[12909];
                
                r_data[12911] <= r_data[12910];
                
                r_data[12912] <= r_data[12911];
                
                r_data[12913] <= r_data[12912];
                
                r_data[12914] <= r_data[12913];
                
                r_data[12915] <= r_data[12914];
                
                r_data[12916] <= r_data[12915];
                
                r_data[12917] <= r_data[12916];
                
                r_data[12918] <= r_data[12917];
                
                r_data[12919] <= r_data[12918];
                
                r_data[12920] <= r_data[12919];
                
                r_data[12921] <= r_data[12920];
                
                r_data[12922] <= r_data[12921];
                
                r_data[12923] <= r_data[12922];
                
                r_data[12924] <= r_data[12923];
                
                r_data[12925] <= r_data[12924];
                
                r_data[12926] <= r_data[12925];
                
                r_data[12927] <= r_data[12926];
                
                r_data[12928] <= r_data[12927];
                
                r_data[12929] <= r_data[12928];
                
                r_data[12930] <= r_data[12929];
                
                r_data[12931] <= r_data[12930];
                
                r_data[12932] <= r_data[12931];
                
                r_data[12933] <= r_data[12932];
                
                r_data[12934] <= r_data[12933];
                
                r_data[12935] <= r_data[12934];
                
                r_data[12936] <= r_data[12935];
                
                r_data[12937] <= r_data[12936];
                
                r_data[12938] <= r_data[12937];
                
                r_data[12939] <= r_data[12938];
                
                r_data[12940] <= r_data[12939];
                
                r_data[12941] <= r_data[12940];
                
                r_data[12942] <= r_data[12941];
                
                r_data[12943] <= r_data[12942];
                
                r_data[12944] <= r_data[12943];
                
                r_data[12945] <= r_data[12944];
                
                r_data[12946] <= r_data[12945];
                
                r_data[12947] <= r_data[12946];
                
                r_data[12948] <= r_data[12947];
                
                r_data[12949] <= r_data[12948];
                
                r_data[12950] <= r_data[12949];
                
                r_data[12951] <= r_data[12950];
                
                r_data[12952] <= r_data[12951];
                
                r_data[12953] <= r_data[12952];
                
                r_data[12954] <= r_data[12953];
                
                r_data[12955] <= r_data[12954];
                
                r_data[12956] <= r_data[12955];
                
                r_data[12957] <= r_data[12956];
                
                r_data[12958] <= r_data[12957];
                
                r_data[12959] <= r_data[12958];
                
                r_data[12960] <= r_data[12959];
                
                r_data[12961] <= r_data[12960];
                
                r_data[12962] <= r_data[12961];
                
                r_data[12963] <= r_data[12962];
                
                r_data[12964] <= r_data[12963];
                
                r_data[12965] <= r_data[12964];
                
                r_data[12966] <= r_data[12965];
                
                r_data[12967] <= r_data[12966];
                
                r_data[12968] <= r_data[12967];
                
                r_data[12969] <= r_data[12968];
                
                r_data[12970] <= r_data[12969];
                
                r_data[12971] <= r_data[12970];
                
                r_data[12972] <= r_data[12971];
                
                r_data[12973] <= r_data[12972];
                
                r_data[12974] <= r_data[12973];
                
                r_data[12975] <= r_data[12974];
                
                r_data[12976] <= r_data[12975];
                
                r_data[12977] <= r_data[12976];
                
                r_data[12978] <= r_data[12977];
                
                r_data[12979] <= r_data[12978];
                
                r_data[12980] <= r_data[12979];
                
                r_data[12981] <= r_data[12980];
                
                r_data[12982] <= r_data[12981];
                
                r_data[12983] <= r_data[12982];
                
                r_data[12984] <= r_data[12983];
                
                r_data[12985] <= r_data[12984];
                
                r_data[12986] <= r_data[12985];
                
                r_data[12987] <= r_data[12986];
                
                r_data[12988] <= r_data[12987];
                
                r_data[12989] <= r_data[12988];
                
                r_data[12990] <= r_data[12989];
                
                r_data[12991] <= r_data[12990];
                
                r_data[12992] <= r_data[12991];
                
                r_data[12993] <= r_data[12992];
                
                r_data[12994] <= r_data[12993];
                
                r_data[12995] <= r_data[12994];
                
                r_data[12996] <= r_data[12995];
                
                r_data[12997] <= r_data[12996];
                
                r_data[12998] <= r_data[12997];
                
                r_data[12999] <= r_data[12998];
                
                r_data[13000] <= r_data[12999];
                
                r_data[13001] <= r_data[13000];
                
                r_data[13002] <= r_data[13001];
                
                r_data[13003] <= r_data[13002];
                
                r_data[13004] <= r_data[13003];
                
                r_data[13005] <= r_data[13004];
                
                r_data[13006] <= r_data[13005];
                
                r_data[13007] <= r_data[13006];
                
                r_data[13008] <= r_data[13007];
                
                r_data[13009] <= r_data[13008];
                
                r_data[13010] <= r_data[13009];
                
                r_data[13011] <= r_data[13010];
                
                r_data[13012] <= r_data[13011];
                
                r_data[13013] <= r_data[13012];
                
                r_data[13014] <= r_data[13013];
                
                r_data[13015] <= r_data[13014];
                
                r_data[13016] <= r_data[13015];
                
                r_data[13017] <= r_data[13016];
                
                r_data[13018] <= r_data[13017];
                
                r_data[13019] <= r_data[13018];
                
                r_data[13020] <= r_data[13019];
                
                r_data[13021] <= r_data[13020];
                
                r_data[13022] <= r_data[13021];
                
                r_data[13023] <= r_data[13022];
                
                r_data[13024] <= r_data[13023];
                
                r_data[13025] <= r_data[13024];
                
                r_data[13026] <= r_data[13025];
                
                r_data[13027] <= r_data[13026];
                
                r_data[13028] <= r_data[13027];
                
                r_data[13029] <= r_data[13028];
                
                r_data[13030] <= r_data[13029];
                
                r_data[13031] <= r_data[13030];
                
                r_data[13032] <= r_data[13031];
                
                r_data[13033] <= r_data[13032];
                
                r_data[13034] <= r_data[13033];
                
                r_data[13035] <= r_data[13034];
                
                r_data[13036] <= r_data[13035];
                
                r_data[13037] <= r_data[13036];
                
                r_data[13038] <= r_data[13037];
                
                r_data[13039] <= r_data[13038];
                
                r_data[13040] <= r_data[13039];
                
                r_data[13041] <= r_data[13040];
                
                r_data[13042] <= r_data[13041];
                
                r_data[13043] <= r_data[13042];
                
                r_data[13044] <= r_data[13043];
                
                r_data[13045] <= r_data[13044];
                
                r_data[13046] <= r_data[13045];
                
                r_data[13047] <= r_data[13046];
                
                r_data[13048] <= r_data[13047];
                
                r_data[13049] <= r_data[13048];
                
                r_data[13050] <= r_data[13049];
                
                r_data[13051] <= r_data[13050];
                
                r_data[13052] <= r_data[13051];
                
                r_data[13053] <= r_data[13052];
                
                r_data[13054] <= r_data[13053];
                
                r_data[13055] <= r_data[13054];
                
                r_data[13056] <= r_data[13055];
                
                r_data[13057] <= r_data[13056];
                
                r_data[13058] <= r_data[13057];
                
                r_data[13059] <= r_data[13058];
                
                r_data[13060] <= r_data[13059];
                
                r_data[13061] <= r_data[13060];
                
                r_data[13062] <= r_data[13061];
                
                r_data[13063] <= r_data[13062];
                
                r_data[13064] <= r_data[13063];
                
                r_data[13065] <= r_data[13064];
                
                r_data[13066] <= r_data[13065];
                
                r_data[13067] <= r_data[13066];
                
                r_data[13068] <= r_data[13067];
                
                r_data[13069] <= r_data[13068];
                
                r_data[13070] <= r_data[13069];
                
                r_data[13071] <= r_data[13070];
                
                r_data[13072] <= r_data[13071];
                
                r_data[13073] <= r_data[13072];
                
                r_data[13074] <= r_data[13073];
                
                r_data[13075] <= r_data[13074];
                
                r_data[13076] <= r_data[13075];
                
                r_data[13077] <= r_data[13076];
                
                r_data[13078] <= r_data[13077];
                
                r_data[13079] <= r_data[13078];
                
                r_data[13080] <= r_data[13079];
                
                r_data[13081] <= r_data[13080];
                
                r_data[13082] <= r_data[13081];
                
                r_data[13083] <= r_data[13082];
                
                r_data[13084] <= r_data[13083];
                
                r_data[13085] <= r_data[13084];
                
                r_data[13086] <= r_data[13085];
                
                r_data[13087] <= r_data[13086];
                
                r_data[13088] <= r_data[13087];
                
                r_data[13089] <= r_data[13088];
                
                r_data[13090] <= r_data[13089];
                
                r_data[13091] <= r_data[13090];
                
                r_data[13092] <= r_data[13091];
                
                r_data[13093] <= r_data[13092];
                
                r_data[13094] <= r_data[13093];
                
                r_data[13095] <= r_data[13094];
                
                r_data[13096] <= r_data[13095];
                
                r_data[13097] <= r_data[13096];
                
                r_data[13098] <= r_data[13097];
                
                r_data[13099] <= r_data[13098];
                
                r_data[13100] <= r_data[13099];
                
                r_data[13101] <= r_data[13100];
                
                r_data[13102] <= r_data[13101];
                
                r_data[13103] <= r_data[13102];
                
                r_data[13104] <= r_data[13103];
                
                r_data[13105] <= r_data[13104];
                
                r_data[13106] <= r_data[13105];
                
                r_data[13107] <= r_data[13106];
                
                r_data[13108] <= r_data[13107];
                
                r_data[13109] <= r_data[13108];
                
                r_data[13110] <= r_data[13109];
                
                r_data[13111] <= r_data[13110];
                
                r_data[13112] <= r_data[13111];
                
                r_data[13113] <= r_data[13112];
                
                r_data[13114] <= r_data[13113];
                
                r_data[13115] <= r_data[13114];
                
                r_data[13116] <= r_data[13115];
                
                r_data[13117] <= r_data[13116];
                
                r_data[13118] <= r_data[13117];
                
                r_data[13119] <= r_data[13118];
                
                r_data[13120] <= r_data[13119];
                
                r_data[13121] <= r_data[13120];
                
                r_data[13122] <= r_data[13121];
                
                r_data[13123] <= r_data[13122];
                
                r_data[13124] <= r_data[13123];
                
                r_data[13125] <= r_data[13124];
                
                r_data[13126] <= r_data[13125];
                
                r_data[13127] <= r_data[13126];
                
                r_data[13128] <= r_data[13127];
                
                r_data[13129] <= r_data[13128];
                
                r_data[13130] <= r_data[13129];
                
                r_data[13131] <= r_data[13130];
                
                r_data[13132] <= r_data[13131];
                
                r_data[13133] <= r_data[13132];
                
                r_data[13134] <= r_data[13133];
                
                r_data[13135] <= r_data[13134];
                
                r_data[13136] <= r_data[13135];
                
                r_data[13137] <= r_data[13136];
                
                r_data[13138] <= r_data[13137];
                
                r_data[13139] <= r_data[13138];
                
                r_data[13140] <= r_data[13139];
                
                r_data[13141] <= r_data[13140];
                
                r_data[13142] <= r_data[13141];
                
                r_data[13143] <= r_data[13142];
                
                r_data[13144] <= r_data[13143];
                
                r_data[13145] <= r_data[13144];
                
                r_data[13146] <= r_data[13145];
                
                r_data[13147] <= r_data[13146];
                
                r_data[13148] <= r_data[13147];
                
                r_data[13149] <= r_data[13148];
                
                r_data[13150] <= r_data[13149];
                
                r_data[13151] <= r_data[13150];
                
                r_data[13152] <= r_data[13151];
                
                r_data[13153] <= r_data[13152];
                
                r_data[13154] <= r_data[13153];
                
                r_data[13155] <= r_data[13154];
                
                r_data[13156] <= r_data[13155];
                
                r_data[13157] <= r_data[13156];
                
                r_data[13158] <= r_data[13157];
                
                r_data[13159] <= r_data[13158];
                
                r_data[13160] <= r_data[13159];
                
                r_data[13161] <= r_data[13160];
                
                r_data[13162] <= r_data[13161];
                
                r_data[13163] <= r_data[13162];
                
                r_data[13164] <= r_data[13163];
                
                r_data[13165] <= r_data[13164];
                
                r_data[13166] <= r_data[13165];
                
                r_data[13167] <= r_data[13166];
                
                r_data[13168] <= r_data[13167];
                
                r_data[13169] <= r_data[13168];
                
                r_data[13170] <= r_data[13169];
                
                r_data[13171] <= r_data[13170];
                
                r_data[13172] <= r_data[13171];
                
                r_data[13173] <= r_data[13172];
                
                r_data[13174] <= r_data[13173];
                
                r_data[13175] <= r_data[13174];
                
                r_data[13176] <= r_data[13175];
                
                r_data[13177] <= r_data[13176];
                
                r_data[13178] <= r_data[13177];
                
                r_data[13179] <= r_data[13178];
                
                r_data[13180] <= r_data[13179];
                
                r_data[13181] <= r_data[13180];
                
                r_data[13182] <= r_data[13181];
                
                r_data[13183] <= r_data[13182];
                
                r_data[13184] <= r_data[13183];
                
                r_data[13185] <= r_data[13184];
                
                r_data[13186] <= r_data[13185];
                
                r_data[13187] <= r_data[13186];
                
                r_data[13188] <= r_data[13187];
                
                r_data[13189] <= r_data[13188];
                
                r_data[13190] <= r_data[13189];
                
                r_data[13191] <= r_data[13190];
                
                r_data[13192] <= r_data[13191];
                
                r_data[13193] <= r_data[13192];
                
                r_data[13194] <= r_data[13193];
                
                r_data[13195] <= r_data[13194];
                
                r_data[13196] <= r_data[13195];
                
                r_data[13197] <= r_data[13196];
                
                r_data[13198] <= r_data[13197];
                
                r_data[13199] <= r_data[13198];
                
                r_data[13200] <= r_data[13199];
                
                r_data[13201] <= r_data[13200];
                
                r_data[13202] <= r_data[13201];
                
                r_data[13203] <= r_data[13202];
                
                r_data[13204] <= r_data[13203];
                
                r_data[13205] <= r_data[13204];
                
                r_data[13206] <= r_data[13205];
                
                r_data[13207] <= r_data[13206];
                
                r_data[13208] <= r_data[13207];
                
                r_data[13209] <= r_data[13208];
                
                r_data[13210] <= r_data[13209];
                
                r_data[13211] <= r_data[13210];
                
                r_data[13212] <= r_data[13211];
                
                r_data[13213] <= r_data[13212];
                
                r_data[13214] <= r_data[13213];
                
                r_data[13215] <= r_data[13214];
                
                r_data[13216] <= r_data[13215];
                
                r_data[13217] <= r_data[13216];
                
                r_data[13218] <= r_data[13217];
                
                r_data[13219] <= r_data[13218];
                
                r_data[13220] <= r_data[13219];
                
                r_data[13221] <= r_data[13220];
                
                r_data[13222] <= r_data[13221];
                
                r_data[13223] <= r_data[13222];
                
                r_data[13224] <= r_data[13223];
                
                r_data[13225] <= r_data[13224];
                
                r_data[13226] <= r_data[13225];
                
                r_data[13227] <= r_data[13226];
                
                r_data[13228] <= r_data[13227];
                
                r_data[13229] <= r_data[13228];
                
                r_data[13230] <= r_data[13229];
                
                r_data[13231] <= r_data[13230];
                
                r_data[13232] <= r_data[13231];
                
                r_data[13233] <= r_data[13232];
                
                r_data[13234] <= r_data[13233];
                
                r_data[13235] <= r_data[13234];
                
                r_data[13236] <= r_data[13235];
                
                r_data[13237] <= r_data[13236];
                
                r_data[13238] <= r_data[13237];
                
                r_data[13239] <= r_data[13238];
                
                r_data[13240] <= r_data[13239];
                
                r_data[13241] <= r_data[13240];
                
                r_data[13242] <= r_data[13241];
                
                r_data[13243] <= r_data[13242];
                
                r_data[13244] <= r_data[13243];
                
                r_data[13245] <= r_data[13244];
                
                r_data[13246] <= r_data[13245];
                
                r_data[13247] <= r_data[13246];
                
                r_data[13248] <= r_data[13247];
                
                r_data[13249] <= r_data[13248];
                
                r_data[13250] <= r_data[13249];
                
                r_data[13251] <= r_data[13250];
                
                r_data[13252] <= r_data[13251];
                
                r_data[13253] <= r_data[13252];
                
                r_data[13254] <= r_data[13253];
                
                r_data[13255] <= r_data[13254];
                
                r_data[13256] <= r_data[13255];
                
                r_data[13257] <= r_data[13256];
                
                r_data[13258] <= r_data[13257];
                
                r_data[13259] <= r_data[13258];
                
                r_data[13260] <= r_data[13259];
                
                r_data[13261] <= r_data[13260];
                
                r_data[13262] <= r_data[13261];
                
                r_data[13263] <= r_data[13262];
                
                r_data[13264] <= r_data[13263];
                
                r_data[13265] <= r_data[13264];
                
                r_data[13266] <= r_data[13265];
                
                r_data[13267] <= r_data[13266];
                
                r_data[13268] <= r_data[13267];
                
                r_data[13269] <= r_data[13268];
                
                r_data[13270] <= r_data[13269];
                
                r_data[13271] <= r_data[13270];
                
                r_data[13272] <= r_data[13271];
                
                r_data[13273] <= r_data[13272];
                
                r_data[13274] <= r_data[13273];
                
                r_data[13275] <= r_data[13274];
                
                r_data[13276] <= r_data[13275];
                
                r_data[13277] <= r_data[13276];
                
                r_data[13278] <= r_data[13277];
                
                r_data[13279] <= r_data[13278];
                
                r_data[13280] <= r_data[13279];
                
                r_data[13281] <= r_data[13280];
                
                r_data[13282] <= r_data[13281];
                
                r_data[13283] <= r_data[13282];
                
                r_data[13284] <= r_data[13283];
                
                r_data[13285] <= r_data[13284];
                
                r_data[13286] <= r_data[13285];
                
                r_data[13287] <= r_data[13286];
                
                r_data[13288] <= r_data[13287];
                
                r_data[13289] <= r_data[13288];
                
                r_data[13290] <= r_data[13289];
                
                r_data[13291] <= r_data[13290];
                
                r_data[13292] <= r_data[13291];
                
                r_data[13293] <= r_data[13292];
                
                r_data[13294] <= r_data[13293];
                
                r_data[13295] <= r_data[13294];
                
                r_data[13296] <= r_data[13295];
                
                r_data[13297] <= r_data[13296];
                
                r_data[13298] <= r_data[13297];
                
                r_data[13299] <= r_data[13298];
                
                r_data[13300] <= r_data[13299];
                
                r_data[13301] <= r_data[13300];
                
                r_data[13302] <= r_data[13301];
                
                r_data[13303] <= r_data[13302];
                
                r_data[13304] <= r_data[13303];
                
                r_data[13305] <= r_data[13304];
                
                r_data[13306] <= r_data[13305];
                
                r_data[13307] <= r_data[13306];
                
                r_data[13308] <= r_data[13307];
                
                r_data[13309] <= r_data[13308];
                
                r_data[13310] <= r_data[13309];
                
                r_data[13311] <= r_data[13310];
                
                r_data[13312] <= r_data[13311];
                
                r_data[13313] <= r_data[13312];
                
                r_data[13314] <= r_data[13313];
                
                r_data[13315] <= r_data[13314];
                
                r_data[13316] <= r_data[13315];
                
                r_data[13317] <= r_data[13316];
                
                r_data[13318] <= r_data[13317];
                
                r_data[13319] <= r_data[13318];
                
                r_data[13320] <= r_data[13319];
                
                r_data[13321] <= r_data[13320];
                
                r_data[13322] <= r_data[13321];
                
                r_data[13323] <= r_data[13322];
                
                r_data[13324] <= r_data[13323];
                
                r_data[13325] <= r_data[13324];
                
                r_data[13326] <= r_data[13325];
                
                r_data[13327] <= r_data[13326];
                
                r_data[13328] <= r_data[13327];
                
                r_data[13329] <= r_data[13328];
                
                r_data[13330] <= r_data[13329];
                
                r_data[13331] <= r_data[13330];
                
                r_data[13332] <= r_data[13331];
                
                r_data[13333] <= r_data[13332];
                
                r_data[13334] <= r_data[13333];
                
                r_data[13335] <= r_data[13334];
                
                r_data[13336] <= r_data[13335];
                
                r_data[13337] <= r_data[13336];
                
                r_data[13338] <= r_data[13337];
                
                r_data[13339] <= r_data[13338];
                
                r_data[13340] <= r_data[13339];
                
                r_data[13341] <= r_data[13340];
                
                r_data[13342] <= r_data[13341];
                
                r_data[13343] <= r_data[13342];
                
                r_data[13344] <= r_data[13343];
                
                r_data[13345] <= r_data[13344];
                
                r_data[13346] <= r_data[13345];
                
                r_data[13347] <= r_data[13346];
                
                r_data[13348] <= r_data[13347];
                
                r_data[13349] <= r_data[13348];
                
                r_data[13350] <= r_data[13349];
                
                r_data[13351] <= r_data[13350];
                
                r_data[13352] <= r_data[13351];
                
                r_data[13353] <= r_data[13352];
                
                r_data[13354] <= r_data[13353];
                
                r_data[13355] <= r_data[13354];
                
                r_data[13356] <= r_data[13355];
                
                r_data[13357] <= r_data[13356];
                
                r_data[13358] <= r_data[13357];
                
                r_data[13359] <= r_data[13358];
                
                r_data[13360] <= r_data[13359];
                
                r_data[13361] <= r_data[13360];
                
                r_data[13362] <= r_data[13361];
                
                r_data[13363] <= r_data[13362];
                
                r_data[13364] <= r_data[13363];
                
                r_data[13365] <= r_data[13364];
                
                r_data[13366] <= r_data[13365];
                
                r_data[13367] <= r_data[13366];
                
                r_data[13368] <= r_data[13367];
                
                r_data[13369] <= r_data[13368];
                
                r_data[13370] <= r_data[13369];
                
                r_data[13371] <= r_data[13370];
                
                r_data[13372] <= r_data[13371];
                
                r_data[13373] <= r_data[13372];
                
                r_data[13374] <= r_data[13373];
                
                r_data[13375] <= r_data[13374];
                
                r_data[13376] <= r_data[13375];
                
                r_data[13377] <= r_data[13376];
                
                r_data[13378] <= r_data[13377];
                
                r_data[13379] <= r_data[13378];
                
                r_data[13380] <= r_data[13379];
                
                r_data[13381] <= r_data[13380];
                
                r_data[13382] <= r_data[13381];
                
                r_data[13383] <= r_data[13382];
                
                r_data[13384] <= r_data[13383];
                
                r_data[13385] <= r_data[13384];
                
                r_data[13386] <= r_data[13385];
                
                r_data[13387] <= r_data[13386];
                
                r_data[13388] <= r_data[13387];
                
                r_data[13389] <= r_data[13388];
                
                r_data[13390] <= r_data[13389];
                
                r_data[13391] <= r_data[13390];
                
                r_data[13392] <= r_data[13391];
                
                r_data[13393] <= r_data[13392];
                
                r_data[13394] <= r_data[13393];
                
                r_data[13395] <= r_data[13394];
                
                r_data[13396] <= r_data[13395];
                
                r_data[13397] <= r_data[13396];
                
                r_data[13398] <= r_data[13397];
                
                r_data[13399] <= r_data[13398];
                
                r_data[13400] <= r_data[13399];
                
                r_data[13401] <= r_data[13400];
                
                r_data[13402] <= r_data[13401];
                
                r_data[13403] <= r_data[13402];
                
                r_data[13404] <= r_data[13403];
                
                r_data[13405] <= r_data[13404];
                
                r_data[13406] <= r_data[13405];
                
                r_data[13407] <= r_data[13406];
                
                r_data[13408] <= r_data[13407];
                
                r_data[13409] <= r_data[13408];
                
                r_data[13410] <= r_data[13409];
                
                r_data[13411] <= r_data[13410];
                
                r_data[13412] <= r_data[13411];
                
                r_data[13413] <= r_data[13412];
                
                r_data[13414] <= r_data[13413];
                
                r_data[13415] <= r_data[13414];
                
                r_data[13416] <= r_data[13415];
                
                r_data[13417] <= r_data[13416];
                
                r_data[13418] <= r_data[13417];
                
                r_data[13419] <= r_data[13418];
                
                r_data[13420] <= r_data[13419];
                
                r_data[13421] <= r_data[13420];
                
                r_data[13422] <= r_data[13421];
                
                r_data[13423] <= r_data[13422];
                
                r_data[13424] <= r_data[13423];
                
                r_data[13425] <= r_data[13424];
                
                r_data[13426] <= r_data[13425];
                
                r_data[13427] <= r_data[13426];
                
                r_data[13428] <= r_data[13427];
                
                r_data[13429] <= r_data[13428];
                
                r_data[13430] <= r_data[13429];
                
                r_data[13431] <= r_data[13430];
                
                r_data[13432] <= r_data[13431];
                
                r_data[13433] <= r_data[13432];
                
                r_data[13434] <= r_data[13433];
                
                r_data[13435] <= r_data[13434];
                
                r_data[13436] <= r_data[13435];
                
                r_data[13437] <= r_data[13436];
                
                r_data[13438] <= r_data[13437];
                
                r_data[13439] <= r_data[13438];
                
                r_data[13440] <= r_data[13439];
                
                r_data[13441] <= r_data[13440];
                
                r_data[13442] <= r_data[13441];
                
                r_data[13443] <= r_data[13442];
                
                r_data[13444] <= r_data[13443];
                
                r_data[13445] <= r_data[13444];
                
                r_data[13446] <= r_data[13445];
                
                r_data[13447] <= r_data[13446];
                
                r_data[13448] <= r_data[13447];
                
                r_data[13449] <= r_data[13448];
                
                r_data[13450] <= r_data[13449];
                
                r_data[13451] <= r_data[13450];
                
                r_data[13452] <= r_data[13451];
                
                r_data[13453] <= r_data[13452];
                
                r_data[13454] <= r_data[13453];
                
                r_data[13455] <= r_data[13454];
                
                r_data[13456] <= r_data[13455];
                
                r_data[13457] <= r_data[13456];
                
                r_data[13458] <= r_data[13457];
                
                r_data[13459] <= r_data[13458];
                
                r_data[13460] <= r_data[13459];
                
                r_data[13461] <= r_data[13460];
                
                r_data[13462] <= r_data[13461];
                
                r_data[13463] <= r_data[13462];
                
                r_data[13464] <= r_data[13463];
                
                r_data[13465] <= r_data[13464];
                
                r_data[13466] <= r_data[13465];
                
                r_data[13467] <= r_data[13466];
                
                r_data[13468] <= r_data[13467];
                
                r_data[13469] <= r_data[13468];
                
                r_data[13470] <= r_data[13469];
                
                r_data[13471] <= r_data[13470];
                
                r_data[13472] <= r_data[13471];
                
                r_data[13473] <= r_data[13472];
                
                r_data[13474] <= r_data[13473];
                
                r_data[13475] <= r_data[13474];
                
                r_data[13476] <= r_data[13475];
                
                r_data[13477] <= r_data[13476];
                
                r_data[13478] <= r_data[13477];
                
                r_data[13479] <= r_data[13478];
                
                r_data[13480] <= r_data[13479];
                
                r_data[13481] <= r_data[13480];
                
                r_data[13482] <= r_data[13481];
                
                r_data[13483] <= r_data[13482];
                
                r_data[13484] <= r_data[13483];
                
                r_data[13485] <= r_data[13484];
                
                r_data[13486] <= r_data[13485];
                
                r_data[13487] <= r_data[13486];
                
                r_data[13488] <= r_data[13487];
                
                r_data[13489] <= r_data[13488];
                
                r_data[13490] <= r_data[13489];
                
                r_data[13491] <= r_data[13490];
                
                r_data[13492] <= r_data[13491];
                
                r_data[13493] <= r_data[13492];
                
                r_data[13494] <= r_data[13493];
                
                r_data[13495] <= r_data[13494];
                
                r_data[13496] <= r_data[13495];
                
                r_data[13497] <= r_data[13496];
                
                r_data[13498] <= r_data[13497];
                
                r_data[13499] <= r_data[13498];
                
                r_data[13500] <= r_data[13499];
                
                r_data[13501] <= r_data[13500];
                
                r_data[13502] <= r_data[13501];
                
                r_data[13503] <= r_data[13502];
                
                r_data[13504] <= r_data[13503];
                
                r_data[13505] <= r_data[13504];
                
                r_data[13506] <= r_data[13505];
                
                r_data[13507] <= r_data[13506];
                
                r_data[13508] <= r_data[13507];
                
                r_data[13509] <= r_data[13508];
                
                r_data[13510] <= r_data[13509];
                
                r_data[13511] <= r_data[13510];
                
                r_data[13512] <= r_data[13511];
                
                r_data[13513] <= r_data[13512];
                
                r_data[13514] <= r_data[13513];
                
                r_data[13515] <= r_data[13514];
                
                r_data[13516] <= r_data[13515];
                
                r_data[13517] <= r_data[13516];
                
                r_data[13518] <= r_data[13517];
                
                r_data[13519] <= r_data[13518];
                
                r_data[13520] <= r_data[13519];
                
                r_data[13521] <= r_data[13520];
                
                r_data[13522] <= r_data[13521];
                
                r_data[13523] <= r_data[13522];
                
                r_data[13524] <= r_data[13523];
                
                r_data[13525] <= r_data[13524];
                
                r_data[13526] <= r_data[13525];
                
                r_data[13527] <= r_data[13526];
                
                r_data[13528] <= r_data[13527];
                
                r_data[13529] <= r_data[13528];
                
                r_data[13530] <= r_data[13529];
                
                r_data[13531] <= r_data[13530];
                
                r_data[13532] <= r_data[13531];
                
                r_data[13533] <= r_data[13532];
                
                r_data[13534] <= r_data[13533];
                
                r_data[13535] <= r_data[13534];
                
                r_data[13536] <= r_data[13535];
                
                r_data[13537] <= r_data[13536];
                
                r_data[13538] <= r_data[13537];
                
                r_data[13539] <= r_data[13538];
                
                r_data[13540] <= r_data[13539];
                
                r_data[13541] <= r_data[13540];
                
                r_data[13542] <= r_data[13541];
                
                r_data[13543] <= r_data[13542];
                
                r_data[13544] <= r_data[13543];
                
                r_data[13545] <= r_data[13544];
                
                r_data[13546] <= r_data[13545];
                
                r_data[13547] <= r_data[13546];
                
                r_data[13548] <= r_data[13547];
                
                r_data[13549] <= r_data[13548];
                
                r_data[13550] <= r_data[13549];
                
                r_data[13551] <= r_data[13550];
                
                r_data[13552] <= r_data[13551];
                
                r_data[13553] <= r_data[13552];
                
                r_data[13554] <= r_data[13553];
                
                r_data[13555] <= r_data[13554];
                
                r_data[13556] <= r_data[13555];
                
                r_data[13557] <= r_data[13556];
                
                r_data[13558] <= r_data[13557];
                
                r_data[13559] <= r_data[13558];
                
                r_data[13560] <= r_data[13559];
                
                r_data[13561] <= r_data[13560];
                
                r_data[13562] <= r_data[13561];
                
                r_data[13563] <= r_data[13562];
                
                r_data[13564] <= r_data[13563];
                
                r_data[13565] <= r_data[13564];
                
                r_data[13566] <= r_data[13565];
                
                r_data[13567] <= r_data[13566];
                
                r_data[13568] <= r_data[13567];
                
                r_data[13569] <= r_data[13568];
                
                r_data[13570] <= r_data[13569];
                
                r_data[13571] <= r_data[13570];
                
                r_data[13572] <= r_data[13571];
                
                r_data[13573] <= r_data[13572];
                
                r_data[13574] <= r_data[13573];
                
                r_data[13575] <= r_data[13574];
                
                r_data[13576] <= r_data[13575];
                
                r_data[13577] <= r_data[13576];
                
                r_data[13578] <= r_data[13577];
                
                r_data[13579] <= r_data[13578];
                
                r_data[13580] <= r_data[13579];
                
                r_data[13581] <= r_data[13580];
                
                r_data[13582] <= r_data[13581];
                
                r_data[13583] <= r_data[13582];
                
                r_data[13584] <= r_data[13583];
                
                r_data[13585] <= r_data[13584];
                
                r_data[13586] <= r_data[13585];
                
                r_data[13587] <= r_data[13586];
                
                r_data[13588] <= r_data[13587];
                
                r_data[13589] <= r_data[13588];
                
                r_data[13590] <= r_data[13589];
                
                r_data[13591] <= r_data[13590];
                
                r_data[13592] <= r_data[13591];
                
                r_data[13593] <= r_data[13592];
                
                r_data[13594] <= r_data[13593];
                
                r_data[13595] <= r_data[13594];
                
                r_data[13596] <= r_data[13595];
                
                r_data[13597] <= r_data[13596];
                
                r_data[13598] <= r_data[13597];
                
                r_data[13599] <= r_data[13598];
                
                r_data[13600] <= r_data[13599];
                
                r_data[13601] <= r_data[13600];
                
                r_data[13602] <= r_data[13601];
                
                r_data[13603] <= r_data[13602];
                
                r_data[13604] <= r_data[13603];
                
                r_data[13605] <= r_data[13604];
                
                r_data[13606] <= r_data[13605];
                
                r_data[13607] <= r_data[13606];
                
                r_data[13608] <= r_data[13607];
                
                r_data[13609] <= r_data[13608];
                
                r_data[13610] <= r_data[13609];
                
                r_data[13611] <= r_data[13610];
                
                r_data[13612] <= r_data[13611];
                
                r_data[13613] <= r_data[13612];
                
                r_data[13614] <= r_data[13613];
                
                r_data[13615] <= r_data[13614];
                
                r_data[13616] <= r_data[13615];
                
                r_data[13617] <= r_data[13616];
                
                r_data[13618] <= r_data[13617];
                
                r_data[13619] <= r_data[13618];
                
                r_data[13620] <= r_data[13619];
                
                r_data[13621] <= r_data[13620];
                
                r_data[13622] <= r_data[13621];
                
                r_data[13623] <= r_data[13622];
                
                r_data[13624] <= r_data[13623];
                
                r_data[13625] <= r_data[13624];
                
                r_data[13626] <= r_data[13625];
                
                r_data[13627] <= r_data[13626];
                
                r_data[13628] <= r_data[13627];
                
                r_data[13629] <= r_data[13628];
                
                r_data[13630] <= r_data[13629];
                
                r_data[13631] <= r_data[13630];
                
                r_data[13632] <= r_data[13631];
                
                r_data[13633] <= r_data[13632];
                
                r_data[13634] <= r_data[13633];
                
                r_data[13635] <= r_data[13634];
                
                r_data[13636] <= r_data[13635];
                
                r_data[13637] <= r_data[13636];
                
                r_data[13638] <= r_data[13637];
                
                r_data[13639] <= r_data[13638];
                
                r_data[13640] <= r_data[13639];
                
                r_data[13641] <= r_data[13640];
                
                r_data[13642] <= r_data[13641];
                
                r_data[13643] <= r_data[13642];
                
                r_data[13644] <= r_data[13643];
                
                r_data[13645] <= r_data[13644];
                
                r_data[13646] <= r_data[13645];
                
                r_data[13647] <= r_data[13646];
                
                r_data[13648] <= r_data[13647];
                
                r_data[13649] <= r_data[13648];
                
                r_data[13650] <= r_data[13649];
                
                r_data[13651] <= r_data[13650];
                
                r_data[13652] <= r_data[13651];
                
                r_data[13653] <= r_data[13652];
                
                r_data[13654] <= r_data[13653];
                
                r_data[13655] <= r_data[13654];
                
                r_data[13656] <= r_data[13655];
                
                r_data[13657] <= r_data[13656];
                
                r_data[13658] <= r_data[13657];
                
                r_data[13659] <= r_data[13658];
                
                r_data[13660] <= r_data[13659];
                
                r_data[13661] <= r_data[13660];
                
                r_data[13662] <= r_data[13661];
                
                r_data[13663] <= r_data[13662];
                
                r_data[13664] <= r_data[13663];
                
                r_data[13665] <= r_data[13664];
                
                r_data[13666] <= r_data[13665];
                
                r_data[13667] <= r_data[13666];
                
                r_data[13668] <= r_data[13667];
                
                r_data[13669] <= r_data[13668];
                
                r_data[13670] <= r_data[13669];
                
                r_data[13671] <= r_data[13670];
                
                r_data[13672] <= r_data[13671];
                
                r_data[13673] <= r_data[13672];
                
                r_data[13674] <= r_data[13673];
                
                r_data[13675] <= r_data[13674];
                
                r_data[13676] <= r_data[13675];
                
                r_data[13677] <= r_data[13676];
                
                r_data[13678] <= r_data[13677];
                
                r_data[13679] <= r_data[13678];
                
                r_data[13680] <= r_data[13679];
                
                r_data[13681] <= r_data[13680];
                
                r_data[13682] <= r_data[13681];
                
                r_data[13683] <= r_data[13682];
                
                r_data[13684] <= r_data[13683];
                
                r_data[13685] <= r_data[13684];
                
                r_data[13686] <= r_data[13685];
                
                r_data[13687] <= r_data[13686];
                
                r_data[13688] <= r_data[13687];
                
                r_data[13689] <= r_data[13688];
                
                r_data[13690] <= r_data[13689];
                
                r_data[13691] <= r_data[13690];
                
                r_data[13692] <= r_data[13691];
                
                r_data[13693] <= r_data[13692];
                
                r_data[13694] <= r_data[13693];
                
                r_data[13695] <= r_data[13694];
                
                r_data[13696] <= r_data[13695];
                
                r_data[13697] <= r_data[13696];
                
                r_data[13698] <= r_data[13697];
                
                r_data[13699] <= r_data[13698];
                
                r_data[13700] <= r_data[13699];
                
                r_data[13701] <= r_data[13700];
                
                r_data[13702] <= r_data[13701];
                
                r_data[13703] <= r_data[13702];
                
                r_data[13704] <= r_data[13703];
                
                r_data[13705] <= r_data[13704];
                
                r_data[13706] <= r_data[13705];
                
                r_data[13707] <= r_data[13706];
                
                r_data[13708] <= r_data[13707];
                
                r_data[13709] <= r_data[13708];
                
                r_data[13710] <= r_data[13709];
                
                r_data[13711] <= r_data[13710];
                
                r_data[13712] <= r_data[13711];
                
                r_data[13713] <= r_data[13712];
                
                r_data[13714] <= r_data[13713];
                
                r_data[13715] <= r_data[13714];
                
                r_data[13716] <= r_data[13715];
                
                r_data[13717] <= r_data[13716];
                
                r_data[13718] <= r_data[13717];
                
                r_data[13719] <= r_data[13718];
                
                r_data[13720] <= r_data[13719];
                
                r_data[13721] <= r_data[13720];
                
                r_data[13722] <= r_data[13721];
                
                r_data[13723] <= r_data[13722];
                
                r_data[13724] <= r_data[13723];
                
                r_data[13725] <= r_data[13724];
                
                r_data[13726] <= r_data[13725];
                
                r_data[13727] <= r_data[13726];
                
                r_data[13728] <= r_data[13727];
                
                r_data[13729] <= r_data[13728];
                
                r_data[13730] <= r_data[13729];
                
                r_data[13731] <= r_data[13730];
                
                r_data[13732] <= r_data[13731];
                
                r_data[13733] <= r_data[13732];
                
                r_data[13734] <= r_data[13733];
                
                r_data[13735] <= r_data[13734];
                
                r_data[13736] <= r_data[13735];
                
                r_data[13737] <= r_data[13736];
                
                r_data[13738] <= r_data[13737];
                
                r_data[13739] <= r_data[13738];
                
                r_data[13740] <= r_data[13739];
                
                r_data[13741] <= r_data[13740];
                
                r_data[13742] <= r_data[13741];
                
                r_data[13743] <= r_data[13742];
                
                r_data[13744] <= r_data[13743];
                
                r_data[13745] <= r_data[13744];
                
                r_data[13746] <= r_data[13745];
                
                r_data[13747] <= r_data[13746];
                
                r_data[13748] <= r_data[13747];
                
                r_data[13749] <= r_data[13748];
                
                r_data[13750] <= r_data[13749];
                
                r_data[13751] <= r_data[13750];
                
                r_data[13752] <= r_data[13751];
                
                r_data[13753] <= r_data[13752];
                
                r_data[13754] <= r_data[13753];
                
                r_data[13755] <= r_data[13754];
                
                r_data[13756] <= r_data[13755];
                
                r_data[13757] <= r_data[13756];
                
                r_data[13758] <= r_data[13757];
                
                r_data[13759] <= r_data[13758];
                
                r_data[13760] <= r_data[13759];
                
                r_data[13761] <= r_data[13760];
                
                r_data[13762] <= r_data[13761];
                
                r_data[13763] <= r_data[13762];
                
                r_data[13764] <= r_data[13763];
                
                r_data[13765] <= r_data[13764];
                
                r_data[13766] <= r_data[13765];
                
                r_data[13767] <= r_data[13766];
                
                r_data[13768] <= r_data[13767];
                
                r_data[13769] <= r_data[13768];
                
                r_data[13770] <= r_data[13769];
                
                r_data[13771] <= r_data[13770];
                
                r_data[13772] <= r_data[13771];
                
                r_data[13773] <= r_data[13772];
                
                r_data[13774] <= r_data[13773];
                
                r_data[13775] <= r_data[13774];
                
                r_data[13776] <= r_data[13775];
                
                r_data[13777] <= r_data[13776];
                
                r_data[13778] <= r_data[13777];
                
                r_data[13779] <= r_data[13778];
                
                r_data[13780] <= r_data[13779];
                
                r_data[13781] <= r_data[13780];
                
                r_data[13782] <= r_data[13781];
                
                r_data[13783] <= r_data[13782];
                
                r_data[13784] <= r_data[13783];
                
                r_data[13785] <= r_data[13784];
                
                r_data[13786] <= r_data[13785];
                
                r_data[13787] <= r_data[13786];
                
                r_data[13788] <= r_data[13787];
                
                r_data[13789] <= r_data[13788];
                
                r_data[13790] <= r_data[13789];
                
                r_data[13791] <= r_data[13790];
                
                r_data[13792] <= r_data[13791];
                
                r_data[13793] <= r_data[13792];
                
                r_data[13794] <= r_data[13793];
                
                r_data[13795] <= r_data[13794];
                
                r_data[13796] <= r_data[13795];
                
                r_data[13797] <= r_data[13796];
                
                r_data[13798] <= r_data[13797];
                
                r_data[13799] <= r_data[13798];
                
                r_data[13800] <= r_data[13799];
                
                r_data[13801] <= r_data[13800];
                
                r_data[13802] <= r_data[13801];
                
                r_data[13803] <= r_data[13802];
                
                r_data[13804] <= r_data[13803];
                
                r_data[13805] <= r_data[13804];
                
                r_data[13806] <= r_data[13805];
                
                r_data[13807] <= r_data[13806];
                
                r_data[13808] <= r_data[13807];
                
                r_data[13809] <= r_data[13808];
                
                r_data[13810] <= r_data[13809];
                
                r_data[13811] <= r_data[13810];
                
                r_data[13812] <= r_data[13811];
                
                r_data[13813] <= r_data[13812];
                
                r_data[13814] <= r_data[13813];
                
                r_data[13815] <= r_data[13814];
                
                r_data[13816] <= r_data[13815];
                
                r_data[13817] <= r_data[13816];
                
                r_data[13818] <= r_data[13817];
                
                r_data[13819] <= r_data[13818];
                
                r_data[13820] <= r_data[13819];
                
                r_data[13821] <= r_data[13820];
                
                r_data[13822] <= r_data[13821];
                
                r_data[13823] <= r_data[13822];
                
                r_data[13824] <= r_data[13823];
                
                r_data[13825] <= r_data[13824];
                
                r_data[13826] <= r_data[13825];
                
                r_data[13827] <= r_data[13826];
                
                r_data[13828] <= r_data[13827];
                
                r_data[13829] <= r_data[13828];
                
                r_data[13830] <= r_data[13829];
                
                r_data[13831] <= r_data[13830];
                
                r_data[13832] <= r_data[13831];
                
                r_data[13833] <= r_data[13832];
                
                r_data[13834] <= r_data[13833];
                
                r_data[13835] <= r_data[13834];
                
                r_data[13836] <= r_data[13835];
                
                r_data[13837] <= r_data[13836];
                
                r_data[13838] <= r_data[13837];
                
                r_data[13839] <= r_data[13838];
                
                r_data[13840] <= r_data[13839];
                
                r_data[13841] <= r_data[13840];
                
                r_data[13842] <= r_data[13841];
                
                r_data[13843] <= r_data[13842];
                
                r_data[13844] <= r_data[13843];
                
                r_data[13845] <= r_data[13844];
                
                r_data[13846] <= r_data[13845];
                
                r_data[13847] <= r_data[13846];
                
                r_data[13848] <= r_data[13847];
                
                r_data[13849] <= r_data[13848];
                
                r_data[13850] <= r_data[13849];
                
                r_data[13851] <= r_data[13850];
                
                r_data[13852] <= r_data[13851];
                
                r_data[13853] <= r_data[13852];
                
                r_data[13854] <= r_data[13853];
                
                r_data[13855] <= r_data[13854];
                
                r_data[13856] <= r_data[13855];
                
                r_data[13857] <= r_data[13856];
                
                r_data[13858] <= r_data[13857];
                
                r_data[13859] <= r_data[13858];
                
                r_data[13860] <= r_data[13859];
                
                r_data[13861] <= r_data[13860];
                
                r_data[13862] <= r_data[13861];
                
                r_data[13863] <= r_data[13862];
                
                r_data[13864] <= r_data[13863];
                
                r_data[13865] <= r_data[13864];
                
                r_data[13866] <= r_data[13865];
                
                r_data[13867] <= r_data[13866];
                
                r_data[13868] <= r_data[13867];
                
                r_data[13869] <= r_data[13868];
                
                r_data[13870] <= r_data[13869];
                
                r_data[13871] <= r_data[13870];
                
                r_data[13872] <= r_data[13871];
                
                r_data[13873] <= r_data[13872];
                
                r_data[13874] <= r_data[13873];
                
                r_data[13875] <= r_data[13874];
                
                r_data[13876] <= r_data[13875];
                
                r_data[13877] <= r_data[13876];
                
                r_data[13878] <= r_data[13877];
                
                r_data[13879] <= r_data[13878];
                
                r_data[13880] <= r_data[13879];
                
                r_data[13881] <= r_data[13880];
                
                r_data[13882] <= r_data[13881];
                
                r_data[13883] <= r_data[13882];
                
                r_data[13884] <= r_data[13883];
                
                r_data[13885] <= r_data[13884];
                
                r_data[13886] <= r_data[13885];
                
                r_data[13887] <= r_data[13886];
                
                r_data[13888] <= r_data[13887];
                
                r_data[13889] <= r_data[13888];
                
                r_data[13890] <= r_data[13889];
                
                r_data[13891] <= r_data[13890];
                
                r_data[13892] <= r_data[13891];
                
                r_data[13893] <= r_data[13892];
                
                r_data[13894] <= r_data[13893];
                
                r_data[13895] <= r_data[13894];
                
                r_data[13896] <= r_data[13895];
                
                r_data[13897] <= r_data[13896];
                
                r_data[13898] <= r_data[13897];
                
                r_data[13899] <= r_data[13898];
                
                r_data[13900] <= r_data[13899];
                
                r_data[13901] <= r_data[13900];
                
                r_data[13902] <= r_data[13901];
                
                r_data[13903] <= r_data[13902];
                
                r_data[13904] <= r_data[13903];
                
                r_data[13905] <= r_data[13904];
                
                r_data[13906] <= r_data[13905];
                
                r_data[13907] <= r_data[13906];
                
                r_data[13908] <= r_data[13907];
                
                r_data[13909] <= r_data[13908];
                
                r_data[13910] <= r_data[13909];
                
                r_data[13911] <= r_data[13910];
                
                r_data[13912] <= r_data[13911];
                
                r_data[13913] <= r_data[13912];
                
                r_data[13914] <= r_data[13913];
                
                r_data[13915] <= r_data[13914];
                
                r_data[13916] <= r_data[13915];
                
                r_data[13917] <= r_data[13916];
                
                r_data[13918] <= r_data[13917];
                
                r_data[13919] <= r_data[13918];
                
                r_data[13920] <= r_data[13919];
                
                r_data[13921] <= r_data[13920];
                
                r_data[13922] <= r_data[13921];
                
                r_data[13923] <= r_data[13922];
                
                r_data[13924] <= r_data[13923];
                
                r_data[13925] <= r_data[13924];
                
                r_data[13926] <= r_data[13925];
                
                r_data[13927] <= r_data[13926];
                
                r_data[13928] <= r_data[13927];
                
                r_data[13929] <= r_data[13928];
                
                r_data[13930] <= r_data[13929];
                
                r_data[13931] <= r_data[13930];
                
                r_data[13932] <= r_data[13931];
                
                r_data[13933] <= r_data[13932];
                
                r_data[13934] <= r_data[13933];
                
                r_data[13935] <= r_data[13934];
                
                r_data[13936] <= r_data[13935];
                
                r_data[13937] <= r_data[13936];
                
                r_data[13938] <= r_data[13937];
                
                r_data[13939] <= r_data[13938];
                
                r_data[13940] <= r_data[13939];
                
                r_data[13941] <= r_data[13940];
                
                r_data[13942] <= r_data[13941];
                
                r_data[13943] <= r_data[13942];
                
                r_data[13944] <= r_data[13943];
                
                r_data[13945] <= r_data[13944];
                
                r_data[13946] <= r_data[13945];
                
                r_data[13947] <= r_data[13946];
                
                r_data[13948] <= r_data[13947];
                
                r_data[13949] <= r_data[13948];
                
                r_data[13950] <= r_data[13949];
                
                r_data[13951] <= r_data[13950];
                
                r_data[13952] <= r_data[13951];
                
                r_data[13953] <= r_data[13952];
                
                r_data[13954] <= r_data[13953];
                
                r_data[13955] <= r_data[13954];
                
                r_data[13956] <= r_data[13955];
                
                r_data[13957] <= r_data[13956];
                
                r_data[13958] <= r_data[13957];
                
                r_data[13959] <= r_data[13958];
                
                r_data[13960] <= r_data[13959];
                
                r_data[13961] <= r_data[13960];
                
                r_data[13962] <= r_data[13961];
                
                r_data[13963] <= r_data[13962];
                
                r_data[13964] <= r_data[13963];
                
                r_data[13965] <= r_data[13964];
                
                r_data[13966] <= r_data[13965];
                
                r_data[13967] <= r_data[13966];
                
                r_data[13968] <= r_data[13967];
                
                r_data[13969] <= r_data[13968];
                
                r_data[13970] <= r_data[13969];
                
                r_data[13971] <= r_data[13970];
                
                r_data[13972] <= r_data[13971];
                
                r_data[13973] <= r_data[13972];
                
                r_data[13974] <= r_data[13973];
                
                r_data[13975] <= r_data[13974];
                
                r_data[13976] <= r_data[13975];
                
                r_data[13977] <= r_data[13976];
                
                r_data[13978] <= r_data[13977];
                
                r_data[13979] <= r_data[13978];
                
                r_data[13980] <= r_data[13979];
                
                r_data[13981] <= r_data[13980];
                
                r_data[13982] <= r_data[13981];
                
                r_data[13983] <= r_data[13982];
                
                r_data[13984] <= r_data[13983];
                
                r_data[13985] <= r_data[13984];
                
                r_data[13986] <= r_data[13985];
                
                r_data[13987] <= r_data[13986];
                
                r_data[13988] <= r_data[13987];
                
                r_data[13989] <= r_data[13988];
                
                r_data[13990] <= r_data[13989];
                
                r_data[13991] <= r_data[13990];
                
                r_data[13992] <= r_data[13991];
                
                r_data[13993] <= r_data[13992];
                
                r_data[13994] <= r_data[13993];
                
                r_data[13995] <= r_data[13994];
                
                r_data[13996] <= r_data[13995];
                
                r_data[13997] <= r_data[13996];
                
                r_data[13998] <= r_data[13997];
                
                r_data[13999] <= r_data[13998];
                
                r_data[14000] <= r_data[13999];
                
                r_data[14001] <= r_data[14000];
                
                r_data[14002] <= r_data[14001];
                
                r_data[14003] <= r_data[14002];
                
                r_data[14004] <= r_data[14003];
                
                r_data[14005] <= r_data[14004];
                
                r_data[14006] <= r_data[14005];
                
                r_data[14007] <= r_data[14006];
                
                r_data[14008] <= r_data[14007];
                
                r_data[14009] <= r_data[14008];
                
                r_data[14010] <= r_data[14009];
                
                r_data[14011] <= r_data[14010];
                
                r_data[14012] <= r_data[14011];
                
                r_data[14013] <= r_data[14012];
                
                r_data[14014] <= r_data[14013];
                
                r_data[14015] <= r_data[14014];
                
                r_data[14016] <= r_data[14015];
                
                r_data[14017] <= r_data[14016];
                
                r_data[14018] <= r_data[14017];
                
                r_data[14019] <= r_data[14018];
                
                r_data[14020] <= r_data[14019];
                
                r_data[14021] <= r_data[14020];
                
                r_data[14022] <= r_data[14021];
                
                r_data[14023] <= r_data[14022];
                
                r_data[14024] <= r_data[14023];
                
                r_data[14025] <= r_data[14024];
                
                r_data[14026] <= r_data[14025];
                
                r_data[14027] <= r_data[14026];
                
                r_data[14028] <= r_data[14027];
                
                r_data[14029] <= r_data[14028];
                
                r_data[14030] <= r_data[14029];
                
                r_data[14031] <= r_data[14030];
                
                r_data[14032] <= r_data[14031];
                
                r_data[14033] <= r_data[14032];
                
                r_data[14034] <= r_data[14033];
                
                r_data[14035] <= r_data[14034];
                
                r_data[14036] <= r_data[14035];
                
                r_data[14037] <= r_data[14036];
                
                r_data[14038] <= r_data[14037];
                
                r_data[14039] <= r_data[14038];
                
                r_data[14040] <= r_data[14039];
                
                r_data[14041] <= r_data[14040];
                
                r_data[14042] <= r_data[14041];
                
                r_data[14043] <= r_data[14042];
                
                r_data[14044] <= r_data[14043];
                
                r_data[14045] <= r_data[14044];
                
                r_data[14046] <= r_data[14045];
                
                r_data[14047] <= r_data[14046];
                
                r_data[14048] <= r_data[14047];
                
                r_data[14049] <= r_data[14048];
                
                r_data[14050] <= r_data[14049];
                
                r_data[14051] <= r_data[14050];
                
                r_data[14052] <= r_data[14051];
                
                r_data[14053] <= r_data[14052];
                
                r_data[14054] <= r_data[14053];
                
                r_data[14055] <= r_data[14054];
                
                r_data[14056] <= r_data[14055];
                
                r_data[14057] <= r_data[14056];
                
                r_data[14058] <= r_data[14057];
                
                r_data[14059] <= r_data[14058];
                
                r_data[14060] <= r_data[14059];
                
                r_data[14061] <= r_data[14060];
                
                r_data[14062] <= r_data[14061];
                
                r_data[14063] <= r_data[14062];
                
                r_data[14064] <= r_data[14063];
                
                r_data[14065] <= r_data[14064];
                
                r_data[14066] <= r_data[14065];
                
                r_data[14067] <= r_data[14066];
                
                r_data[14068] <= r_data[14067];
                
                r_data[14069] <= r_data[14068];
                
                r_data[14070] <= r_data[14069];
                
                r_data[14071] <= r_data[14070];
                
                r_data[14072] <= r_data[14071];
                
                r_data[14073] <= r_data[14072];
                
                r_data[14074] <= r_data[14073];
                
                r_data[14075] <= r_data[14074];
                
                r_data[14076] <= r_data[14075];
                
                r_data[14077] <= r_data[14076];
                
                r_data[14078] <= r_data[14077];
                
                r_data[14079] <= r_data[14078];
                
                r_data[14080] <= r_data[14079];
                
                r_data[14081] <= r_data[14080];
                
                r_data[14082] <= r_data[14081];
                
                r_data[14083] <= r_data[14082];
                
                r_data[14084] <= r_data[14083];
                
                r_data[14085] <= r_data[14084];
                
                r_data[14086] <= r_data[14085];
                
                r_data[14087] <= r_data[14086];
                
                r_data[14088] <= r_data[14087];
                
                r_data[14089] <= r_data[14088];
                
                r_data[14090] <= r_data[14089];
                
                r_data[14091] <= r_data[14090];
                
                r_data[14092] <= r_data[14091];
                
                r_data[14093] <= r_data[14092];
                
                r_data[14094] <= r_data[14093];
                
                r_data[14095] <= r_data[14094];
                
                r_data[14096] <= r_data[14095];
                
                r_data[14097] <= r_data[14096];
                
                r_data[14098] <= r_data[14097];
                
                r_data[14099] <= r_data[14098];
                
                r_data[14100] <= r_data[14099];
                
                r_data[14101] <= r_data[14100];
                
                r_data[14102] <= r_data[14101];
                
                r_data[14103] <= r_data[14102];
                
                r_data[14104] <= r_data[14103];
                
                r_data[14105] <= r_data[14104];
                
                r_data[14106] <= r_data[14105];
                
                r_data[14107] <= r_data[14106];
                
                r_data[14108] <= r_data[14107];
                
                r_data[14109] <= r_data[14108];
                
                r_data[14110] <= r_data[14109];
                
                r_data[14111] <= r_data[14110];
                
                r_data[14112] <= r_data[14111];
                
                r_data[14113] <= r_data[14112];
                
                r_data[14114] <= r_data[14113];
                
                r_data[14115] <= r_data[14114];
                
                r_data[14116] <= r_data[14115];
                
                r_data[14117] <= r_data[14116];
                
                r_data[14118] <= r_data[14117];
                
                r_data[14119] <= r_data[14118];
                
                r_data[14120] <= r_data[14119];
                
                r_data[14121] <= r_data[14120];
                
                r_data[14122] <= r_data[14121];
                
                r_data[14123] <= r_data[14122];
                
                r_data[14124] <= r_data[14123];
                
                r_data[14125] <= r_data[14124];
                
                r_data[14126] <= r_data[14125];
                
                r_data[14127] <= r_data[14126];
                
                r_data[14128] <= r_data[14127];
                
                r_data[14129] <= r_data[14128];
                
                r_data[14130] <= r_data[14129];
                
                r_data[14131] <= r_data[14130];
                
                r_data[14132] <= r_data[14131];
                
                r_data[14133] <= r_data[14132];
                
                r_data[14134] <= r_data[14133];
                
                r_data[14135] <= r_data[14134];
                
                r_data[14136] <= r_data[14135];
                
                r_data[14137] <= r_data[14136];
                
                r_data[14138] <= r_data[14137];
                
                r_data[14139] <= r_data[14138];
                
                r_data[14140] <= r_data[14139];
                
                r_data[14141] <= r_data[14140];
                
                r_data[14142] <= r_data[14141];
                
                r_data[14143] <= r_data[14142];
                
                r_data[14144] <= r_data[14143];
                
                r_data[14145] <= r_data[14144];
                
                r_data[14146] <= r_data[14145];
                
                r_data[14147] <= r_data[14146];
                
                r_data[14148] <= r_data[14147];
                
                r_data[14149] <= r_data[14148];
                
                r_data[14150] <= r_data[14149];
                
                r_data[14151] <= r_data[14150];
                
                r_data[14152] <= r_data[14151];
                
                r_data[14153] <= r_data[14152];
                
                r_data[14154] <= r_data[14153];
                
                r_data[14155] <= r_data[14154];
                
                r_data[14156] <= r_data[14155];
                
                r_data[14157] <= r_data[14156];
                
                r_data[14158] <= r_data[14157];
                
                r_data[14159] <= r_data[14158];
                
                r_data[14160] <= r_data[14159];
                
                r_data[14161] <= r_data[14160];
                
                r_data[14162] <= r_data[14161];
                
                r_data[14163] <= r_data[14162];
                
                r_data[14164] <= r_data[14163];
                
                r_data[14165] <= r_data[14164];
                
                r_data[14166] <= r_data[14165];
                
                r_data[14167] <= r_data[14166];
                
                r_data[14168] <= r_data[14167];
                
                r_data[14169] <= r_data[14168];
                
                r_data[14170] <= r_data[14169];
                
                r_data[14171] <= r_data[14170];
                
                r_data[14172] <= r_data[14171];
                
                r_data[14173] <= r_data[14172];
                
                r_data[14174] <= r_data[14173];
                
                r_data[14175] <= r_data[14174];
                
                r_data[14176] <= r_data[14175];
                
                r_data[14177] <= r_data[14176];
                
                r_data[14178] <= r_data[14177];
                
                r_data[14179] <= r_data[14178];
                
                r_data[14180] <= r_data[14179];
                
                r_data[14181] <= r_data[14180];
                
                r_data[14182] <= r_data[14181];
                
                r_data[14183] <= r_data[14182];
                
                r_data[14184] <= r_data[14183];
                
                r_data[14185] <= r_data[14184];
                
                r_data[14186] <= r_data[14185];
                
                r_data[14187] <= r_data[14186];
                
                r_data[14188] <= r_data[14187];
                
                r_data[14189] <= r_data[14188];
                
                r_data[14190] <= r_data[14189];
                
                r_data[14191] <= r_data[14190];
                
                r_data[14192] <= r_data[14191];
                
                r_data[14193] <= r_data[14192];
                
                r_data[14194] <= r_data[14193];
                
                r_data[14195] <= r_data[14194];
                
                r_data[14196] <= r_data[14195];
                
                r_data[14197] <= r_data[14196];
                
                r_data[14198] <= r_data[14197];
                
                r_data[14199] <= r_data[14198];
                
                r_data[14200] <= r_data[14199];
                
                r_data[14201] <= r_data[14200];
                
                r_data[14202] <= r_data[14201];
                
                r_data[14203] <= r_data[14202];
                
                r_data[14204] <= r_data[14203];
                
                r_data[14205] <= r_data[14204];
                
                r_data[14206] <= r_data[14205];
                
                r_data[14207] <= r_data[14206];
                
                r_data[14208] <= r_data[14207];
                
                r_data[14209] <= r_data[14208];
                
                r_data[14210] <= r_data[14209];
                
                r_data[14211] <= r_data[14210];
                
                r_data[14212] <= r_data[14211];
                
                r_data[14213] <= r_data[14212];
                
                r_data[14214] <= r_data[14213];
                
                r_data[14215] <= r_data[14214];
                
                r_data[14216] <= r_data[14215];
                
                r_data[14217] <= r_data[14216];
                
                r_data[14218] <= r_data[14217];
                
                r_data[14219] <= r_data[14218];
                
                r_data[14220] <= r_data[14219];
                
                r_data[14221] <= r_data[14220];
                
                r_data[14222] <= r_data[14221];
                
                r_data[14223] <= r_data[14222];
                
                r_data[14224] <= r_data[14223];
                
                r_data[14225] <= r_data[14224];
                
                r_data[14226] <= r_data[14225];
                
                r_data[14227] <= r_data[14226];
                
                r_data[14228] <= r_data[14227];
                
                r_data[14229] <= r_data[14228];
                
                r_data[14230] <= r_data[14229];
                
                r_data[14231] <= r_data[14230];
                
                r_data[14232] <= r_data[14231];
                
                r_data[14233] <= r_data[14232];
                
                r_data[14234] <= r_data[14233];
                
                r_data[14235] <= r_data[14234];
                
                r_data[14236] <= r_data[14235];
                
                r_data[14237] <= r_data[14236];
                
                r_data[14238] <= r_data[14237];
                
                r_data[14239] <= r_data[14238];
                
                r_data[14240] <= r_data[14239];
                
                r_data[14241] <= r_data[14240];
                
                r_data[14242] <= r_data[14241];
                
                r_data[14243] <= r_data[14242];
                
                r_data[14244] <= r_data[14243];
                
                r_data[14245] <= r_data[14244];
                
                r_data[14246] <= r_data[14245];
                
                r_data[14247] <= r_data[14246];
                
                r_data[14248] <= r_data[14247];
                
                r_data[14249] <= r_data[14248];
                
                r_data[14250] <= r_data[14249];
                
                r_data[14251] <= r_data[14250];
                
                r_data[14252] <= r_data[14251];
                
                r_data[14253] <= r_data[14252];
                
                r_data[14254] <= r_data[14253];
                
                r_data[14255] <= r_data[14254];
                
                r_data[14256] <= r_data[14255];
                
                r_data[14257] <= r_data[14256];
                
                r_data[14258] <= r_data[14257];
                
                r_data[14259] <= r_data[14258];
                
                r_data[14260] <= r_data[14259];
                
                r_data[14261] <= r_data[14260];
                
                r_data[14262] <= r_data[14261];
                
                r_data[14263] <= r_data[14262];
                
                r_data[14264] <= r_data[14263];
                
                r_data[14265] <= r_data[14264];
                
                r_data[14266] <= r_data[14265];
                
                r_data[14267] <= r_data[14266];
                
                r_data[14268] <= r_data[14267];
                
                r_data[14269] <= r_data[14268];
                
                r_data[14270] <= r_data[14269];
                
                r_data[14271] <= r_data[14270];
                
                r_data[14272] <= r_data[14271];
                
                r_data[14273] <= r_data[14272];
                
                r_data[14274] <= r_data[14273];
                
                r_data[14275] <= r_data[14274];
                
                r_data[14276] <= r_data[14275];
                
                r_data[14277] <= r_data[14276];
                
                r_data[14278] <= r_data[14277];
                
                r_data[14279] <= r_data[14278];
                
                r_data[14280] <= r_data[14279];
                
                r_data[14281] <= r_data[14280];
                
                r_data[14282] <= r_data[14281];
                
                r_data[14283] <= r_data[14282];
                
                r_data[14284] <= r_data[14283];
                
                r_data[14285] <= r_data[14284];
                
                r_data[14286] <= r_data[14285];
                
                r_data[14287] <= r_data[14286];
                
                r_data[14288] <= r_data[14287];
                
                r_data[14289] <= r_data[14288];
                
                r_data[14290] <= r_data[14289];
                
                r_data[14291] <= r_data[14290];
                
                r_data[14292] <= r_data[14291];
                
                r_data[14293] <= r_data[14292];
                
                r_data[14294] <= r_data[14293];
                
                r_data[14295] <= r_data[14294];
                
                r_data[14296] <= r_data[14295];
                
                r_data[14297] <= r_data[14296];
                
                r_data[14298] <= r_data[14297];
                
                r_data[14299] <= r_data[14298];
                
                r_data[14300] <= r_data[14299];
                
                r_data[14301] <= r_data[14300];
                
                r_data[14302] <= r_data[14301];
                
                r_data[14303] <= r_data[14302];
                
                r_data[14304] <= r_data[14303];
                
                r_data[14305] <= r_data[14304];
                
                r_data[14306] <= r_data[14305];
                
                r_data[14307] <= r_data[14306];
                
                r_data[14308] <= r_data[14307];
                
                r_data[14309] <= r_data[14308];
                
                r_data[14310] <= r_data[14309];
                
                r_data[14311] <= r_data[14310];
                
                r_data[14312] <= r_data[14311];
                
                r_data[14313] <= r_data[14312];
                
                r_data[14314] <= r_data[14313];
                
                r_data[14315] <= r_data[14314];
                
                r_data[14316] <= r_data[14315];
                
                r_data[14317] <= r_data[14316];
                
                r_data[14318] <= r_data[14317];
                
                r_data[14319] <= r_data[14318];
                
                r_data[14320] <= r_data[14319];
                
                r_data[14321] <= r_data[14320];
                
                r_data[14322] <= r_data[14321];
                
                r_data[14323] <= r_data[14322];
                
                r_data[14324] <= r_data[14323];
                
                r_data[14325] <= r_data[14324];
                
                r_data[14326] <= r_data[14325];
                
                r_data[14327] <= r_data[14326];
                
                r_data[14328] <= r_data[14327];
                
                r_data[14329] <= r_data[14328];
                
                r_data[14330] <= r_data[14329];
                
                r_data[14331] <= r_data[14330];
                
                r_data[14332] <= r_data[14331];
                
                r_data[14333] <= r_data[14332];
                
                r_data[14334] <= r_data[14333];
                
                r_data[14335] <= r_data[14334];
                
                r_data[14336] <= r_data[14335];
                
                r_data[14337] <= r_data[14336];
                
                r_data[14338] <= r_data[14337];
                
                r_data[14339] <= r_data[14338];
                
                r_data[14340] <= r_data[14339];
                
                r_data[14341] <= r_data[14340];
                
                r_data[14342] <= r_data[14341];
                
                r_data[14343] <= r_data[14342];
                
                r_data[14344] <= r_data[14343];
                
                r_data[14345] <= r_data[14344];
                
                r_data[14346] <= r_data[14345];
                
                r_data[14347] <= r_data[14346];
                
                r_data[14348] <= r_data[14347];
                
                r_data[14349] <= r_data[14348];
                
                r_data[14350] <= r_data[14349];
                
                r_data[14351] <= r_data[14350];
                
                r_data[14352] <= r_data[14351];
                
                r_data[14353] <= r_data[14352];
                
                r_data[14354] <= r_data[14353];
                
                r_data[14355] <= r_data[14354];
                
                r_data[14356] <= r_data[14355];
                
                r_data[14357] <= r_data[14356];
                
                r_data[14358] <= r_data[14357];
                
                r_data[14359] <= r_data[14358];
                
                r_data[14360] <= r_data[14359];
                
                r_data[14361] <= r_data[14360];
                
                r_data[14362] <= r_data[14361];
                
                r_data[14363] <= r_data[14362];
                
                r_data[14364] <= r_data[14363];
                
                r_data[14365] <= r_data[14364];
                
                r_data[14366] <= r_data[14365];
                
                r_data[14367] <= r_data[14366];
                
                r_data[14368] <= r_data[14367];
                
                r_data[14369] <= r_data[14368];
                
                r_data[14370] <= r_data[14369];
                
                r_data[14371] <= r_data[14370];
                
                r_data[14372] <= r_data[14371];
                
                r_data[14373] <= r_data[14372];
                
                r_data[14374] <= r_data[14373];
                
                r_data[14375] <= r_data[14374];
                
                r_data[14376] <= r_data[14375];
                
                r_data[14377] <= r_data[14376];
                
                r_data[14378] <= r_data[14377];
                
                r_data[14379] <= r_data[14378];
                
                r_data[14380] <= r_data[14379];
                
                r_data[14381] <= r_data[14380];
                
                r_data[14382] <= r_data[14381];
                
                r_data[14383] <= r_data[14382];
                
                r_data[14384] <= r_data[14383];
                
                r_data[14385] <= r_data[14384];
                
                r_data[14386] <= r_data[14385];
                
                r_data[14387] <= r_data[14386];
                
                r_data[14388] <= r_data[14387];
                
                r_data[14389] <= r_data[14388];
                
                r_data[14390] <= r_data[14389];
                
                r_data[14391] <= r_data[14390];
                
                r_data[14392] <= r_data[14391];
                
                r_data[14393] <= r_data[14392];
                
                r_data[14394] <= r_data[14393];
                
                r_data[14395] <= r_data[14394];
                
                r_data[14396] <= r_data[14395];
                
                r_data[14397] <= r_data[14396];
                
                r_data[14398] <= r_data[14397];
                
                r_data[14399] <= r_data[14398];
                
                r_data[14400] <= r_data[14399];
                
                r_data[14401] <= r_data[14400];
                
                r_data[14402] <= r_data[14401];
                
                r_data[14403] <= r_data[14402];
                
                r_data[14404] <= r_data[14403];
                
                r_data[14405] <= r_data[14404];
                
                r_data[14406] <= r_data[14405];
                
                r_data[14407] <= r_data[14406];
                
                r_data[14408] <= r_data[14407];
                
                r_data[14409] <= r_data[14408];
                
                r_data[14410] <= r_data[14409];
                
                r_data[14411] <= r_data[14410];
                
                r_data[14412] <= r_data[14411];
                
                r_data[14413] <= r_data[14412];
                
                r_data[14414] <= r_data[14413];
                
                r_data[14415] <= r_data[14414];
                
                r_data[14416] <= r_data[14415];
                
                r_data[14417] <= r_data[14416];
                
                r_data[14418] <= r_data[14417];
                
                r_data[14419] <= r_data[14418];
                
                r_data[14420] <= r_data[14419];
                
                r_data[14421] <= r_data[14420];
                
                r_data[14422] <= r_data[14421];
                
                r_data[14423] <= r_data[14422];
                
                r_data[14424] <= r_data[14423];
                
                r_data[14425] <= r_data[14424];
                
                r_data[14426] <= r_data[14425];
                
                r_data[14427] <= r_data[14426];
                
                r_data[14428] <= r_data[14427];
                
                r_data[14429] <= r_data[14428];
                
                r_data[14430] <= r_data[14429];
                
                r_data[14431] <= r_data[14430];
                
                r_data[14432] <= r_data[14431];
                
                r_data[14433] <= r_data[14432];
                
                r_data[14434] <= r_data[14433];
                
                r_data[14435] <= r_data[14434];
                
                r_data[14436] <= r_data[14435];
                
                r_data[14437] <= r_data[14436];
                
                r_data[14438] <= r_data[14437];
                
                r_data[14439] <= r_data[14438];
                
                r_data[14440] <= r_data[14439];
                
                r_data[14441] <= r_data[14440];
                
                r_data[14442] <= r_data[14441];
                
                r_data[14443] <= r_data[14442];
                
                r_data[14444] <= r_data[14443];
                
                r_data[14445] <= r_data[14444];
                
                r_data[14446] <= r_data[14445];
                
                r_data[14447] <= r_data[14446];
                
                r_data[14448] <= r_data[14447];
                
                r_data[14449] <= r_data[14448];
                
                r_data[14450] <= r_data[14449];
                
                r_data[14451] <= r_data[14450];
                
                r_data[14452] <= r_data[14451];
                
                r_data[14453] <= r_data[14452];
                
                r_data[14454] <= r_data[14453];
                
                r_data[14455] <= r_data[14454];
                
                r_data[14456] <= r_data[14455];
                
                r_data[14457] <= r_data[14456];
                
                r_data[14458] <= r_data[14457];
                
                r_data[14459] <= r_data[14458];
                
                r_data[14460] <= r_data[14459];
                
                r_data[14461] <= r_data[14460];
                
                r_data[14462] <= r_data[14461];
                
                r_data[14463] <= r_data[14462];
                
                r_data[14464] <= r_data[14463];
                
                r_data[14465] <= r_data[14464];
                
                r_data[14466] <= r_data[14465];
                
                r_data[14467] <= r_data[14466];
                
                r_data[14468] <= r_data[14467];
                
                r_data[14469] <= r_data[14468];
                
                r_data[14470] <= r_data[14469];
                
                r_data[14471] <= r_data[14470];
                
                r_data[14472] <= r_data[14471];
                
                r_data[14473] <= r_data[14472];
                
                r_data[14474] <= r_data[14473];
                
                r_data[14475] <= r_data[14474];
                
                r_data[14476] <= r_data[14475];
                
                r_data[14477] <= r_data[14476];
                
                r_data[14478] <= r_data[14477];
                
                r_data[14479] <= r_data[14478];
                
                r_data[14480] <= r_data[14479];
                
                r_data[14481] <= r_data[14480];
                
                r_data[14482] <= r_data[14481];
                
                r_data[14483] <= r_data[14482];
                
                r_data[14484] <= r_data[14483];
                
                r_data[14485] <= r_data[14484];
                
                r_data[14486] <= r_data[14485];
                
                r_data[14487] <= r_data[14486];
                
                r_data[14488] <= r_data[14487];
                
                r_data[14489] <= r_data[14488];
                
                r_data[14490] <= r_data[14489];
                
                r_data[14491] <= r_data[14490];
                
                r_data[14492] <= r_data[14491];
                
                r_data[14493] <= r_data[14492];
                
                r_data[14494] <= r_data[14493];
                
                r_data[14495] <= r_data[14494];
                
                r_data[14496] <= r_data[14495];
                
                r_data[14497] <= r_data[14496];
                
                r_data[14498] <= r_data[14497];
                
                r_data[14499] <= r_data[14498];
                
                r_data[14500] <= r_data[14499];
                
                r_data[14501] <= r_data[14500];
                
                r_data[14502] <= r_data[14501];
                
                r_data[14503] <= r_data[14502];
                
                r_data[14504] <= r_data[14503];
                
                r_data[14505] <= r_data[14504];
                
                r_data[14506] <= r_data[14505];
                
                r_data[14507] <= r_data[14506];
                
                r_data[14508] <= r_data[14507];
                
                r_data[14509] <= r_data[14508];
                
                r_data[14510] <= r_data[14509];
                
                r_data[14511] <= r_data[14510];
                
                r_data[14512] <= r_data[14511];
                
                r_data[14513] <= r_data[14512];
                
                r_data[14514] <= r_data[14513];
                
                r_data[14515] <= r_data[14514];
                
                r_data[14516] <= r_data[14515];
                
                r_data[14517] <= r_data[14516];
                
                r_data[14518] <= r_data[14517];
                
                r_data[14519] <= r_data[14518];
                
                r_data[14520] <= r_data[14519];
                
                r_data[14521] <= r_data[14520];
                
                r_data[14522] <= r_data[14521];
                
                r_data[14523] <= r_data[14522];
                
                r_data[14524] <= r_data[14523];
                
                r_data[14525] <= r_data[14524];
                
                r_data[14526] <= r_data[14525];
                
                r_data[14527] <= r_data[14526];
                
                r_data[14528] <= r_data[14527];
                
                r_data[14529] <= r_data[14528];
                
                r_data[14530] <= r_data[14529];
                
                r_data[14531] <= r_data[14530];
                
                r_data[14532] <= r_data[14531];
                
                r_data[14533] <= r_data[14532];
                
                r_data[14534] <= r_data[14533];
                
                r_data[14535] <= r_data[14534];
                
                r_data[14536] <= r_data[14535];
                
                r_data[14537] <= r_data[14536];
                
                r_data[14538] <= r_data[14537];
                
                r_data[14539] <= r_data[14538];
                
                r_data[14540] <= r_data[14539];
                
                r_data[14541] <= r_data[14540];
                
                r_data[14542] <= r_data[14541];
                
                r_data[14543] <= r_data[14542];
                
                r_data[14544] <= r_data[14543];
                
                r_data[14545] <= r_data[14544];
                
                r_data[14546] <= r_data[14545];
                
                r_data[14547] <= r_data[14546];
                
                r_data[14548] <= r_data[14547];
                
                r_data[14549] <= r_data[14548];
                
                r_data[14550] <= r_data[14549];
                
                r_data[14551] <= r_data[14550];
                
                r_data[14552] <= r_data[14551];
                
                r_data[14553] <= r_data[14552];
                
                r_data[14554] <= r_data[14553];
                
                r_data[14555] <= r_data[14554];
                
                r_data[14556] <= r_data[14555];
                
                r_data[14557] <= r_data[14556];
                
                r_data[14558] <= r_data[14557];
                
                r_data[14559] <= r_data[14558];
                
                r_data[14560] <= r_data[14559];
                
                r_data[14561] <= r_data[14560];
                
                r_data[14562] <= r_data[14561];
                
                r_data[14563] <= r_data[14562];
                
                r_data[14564] <= r_data[14563];
                
                r_data[14565] <= r_data[14564];
                
                r_data[14566] <= r_data[14565];
                
                r_data[14567] <= r_data[14566];
                
                r_data[14568] <= r_data[14567];
                
                r_data[14569] <= r_data[14568];
                
                r_data[14570] <= r_data[14569];
                
                r_data[14571] <= r_data[14570];
                
                r_data[14572] <= r_data[14571];
                
                r_data[14573] <= r_data[14572];
                
                r_data[14574] <= r_data[14573];
                
                r_data[14575] <= r_data[14574];
                
                r_data[14576] <= r_data[14575];
                
                r_data[14577] <= r_data[14576];
                
                r_data[14578] <= r_data[14577];
                
                r_data[14579] <= r_data[14578];
                
                r_data[14580] <= r_data[14579];
                
                r_data[14581] <= r_data[14580];
                
                r_data[14582] <= r_data[14581];
                
                r_data[14583] <= r_data[14582];
                
                r_data[14584] <= r_data[14583];
                
                r_data[14585] <= r_data[14584];
                
                r_data[14586] <= r_data[14585];
                
                r_data[14587] <= r_data[14586];
                
                r_data[14588] <= r_data[14587];
                
                r_data[14589] <= r_data[14588];
                
                r_data[14590] <= r_data[14589];
                
                r_data[14591] <= r_data[14590];
                
                r_data[14592] <= r_data[14591];
                
                r_data[14593] <= r_data[14592];
                
                r_data[14594] <= r_data[14593];
                
                r_data[14595] <= r_data[14594];
                
                r_data[14596] <= r_data[14595];
                
                r_data[14597] <= r_data[14596];
                
                r_data[14598] <= r_data[14597];
                
                r_data[14599] <= r_data[14598];
                
                r_data[14600] <= r_data[14599];
                
                r_data[14601] <= r_data[14600];
                
                r_data[14602] <= r_data[14601];
                
                r_data[14603] <= r_data[14602];
                
                r_data[14604] <= r_data[14603];
                
                r_data[14605] <= r_data[14604];
                
                r_data[14606] <= r_data[14605];
                
                r_data[14607] <= r_data[14606];
                
                r_data[14608] <= r_data[14607];
                
                r_data[14609] <= r_data[14608];
                
                r_data[14610] <= r_data[14609];
                
                r_data[14611] <= r_data[14610];
                
                r_data[14612] <= r_data[14611];
                
                r_data[14613] <= r_data[14612];
                
                r_data[14614] <= r_data[14613];
                
                r_data[14615] <= r_data[14614];
                
                r_data[14616] <= r_data[14615];
                
                r_data[14617] <= r_data[14616];
                
                r_data[14618] <= r_data[14617];
                
                r_data[14619] <= r_data[14618];
                
                r_data[14620] <= r_data[14619];
                
                r_data[14621] <= r_data[14620];
                
                r_data[14622] <= r_data[14621];
                
                r_data[14623] <= r_data[14622];
                
                r_data[14624] <= r_data[14623];
                
                r_data[14625] <= r_data[14624];
                
                r_data[14626] <= r_data[14625];
                
                r_data[14627] <= r_data[14626];
                
                r_data[14628] <= r_data[14627];
                
                r_data[14629] <= r_data[14628];
                
                r_data[14630] <= r_data[14629];
                
                r_data[14631] <= r_data[14630];
                
                r_data[14632] <= r_data[14631];
                
                r_data[14633] <= r_data[14632];
                
                r_data[14634] <= r_data[14633];
                
                r_data[14635] <= r_data[14634];
                
                r_data[14636] <= r_data[14635];
                
                r_data[14637] <= r_data[14636];
                
                r_data[14638] <= r_data[14637];
                
                r_data[14639] <= r_data[14638];
                
                r_data[14640] <= r_data[14639];
                
                r_data[14641] <= r_data[14640];
                
                r_data[14642] <= r_data[14641];
                
                r_data[14643] <= r_data[14642];
                
                r_data[14644] <= r_data[14643];
                
                r_data[14645] <= r_data[14644];
                
                r_data[14646] <= r_data[14645];
                
                r_data[14647] <= r_data[14646];
                
                r_data[14648] <= r_data[14647];
                
                r_data[14649] <= r_data[14648];
                
                r_data[14650] <= r_data[14649];
                
                r_data[14651] <= r_data[14650];
                
                r_data[14652] <= r_data[14651];
                
                r_data[14653] <= r_data[14652];
                
                r_data[14654] <= r_data[14653];
                
                r_data[14655] <= r_data[14654];
                
                r_data[14656] <= r_data[14655];
                
                r_data[14657] <= r_data[14656];
                
                r_data[14658] <= r_data[14657];
                
                r_data[14659] <= r_data[14658];
                
                r_data[14660] <= r_data[14659];
                
                r_data[14661] <= r_data[14660];
                
                r_data[14662] <= r_data[14661];
                
                r_data[14663] <= r_data[14662];
                
                r_data[14664] <= r_data[14663];
                
                r_data[14665] <= r_data[14664];
                
                r_data[14666] <= r_data[14665];
                
                r_data[14667] <= r_data[14666];
                
                r_data[14668] <= r_data[14667];
                
                r_data[14669] <= r_data[14668];
                
                r_data[14670] <= r_data[14669];
                
                r_data[14671] <= r_data[14670];
                
                r_data[14672] <= r_data[14671];
                
                r_data[14673] <= r_data[14672];
                
                r_data[14674] <= r_data[14673];
                
                r_data[14675] <= r_data[14674];
                
                r_data[14676] <= r_data[14675];
                
                r_data[14677] <= r_data[14676];
                
                r_data[14678] <= r_data[14677];
                
                r_data[14679] <= r_data[14678];
                
                r_data[14680] <= r_data[14679];
                
                r_data[14681] <= r_data[14680];
                
                r_data[14682] <= r_data[14681];
                
                r_data[14683] <= r_data[14682];
                
                r_data[14684] <= r_data[14683];
                
                r_data[14685] <= r_data[14684];
                
                r_data[14686] <= r_data[14685];
                
                r_data[14687] <= r_data[14686];
                
                r_data[14688] <= r_data[14687];
                
                r_data[14689] <= r_data[14688];
                
                r_data[14690] <= r_data[14689];
                
                r_data[14691] <= r_data[14690];
                
                r_data[14692] <= r_data[14691];
                
                r_data[14693] <= r_data[14692];
                
                r_data[14694] <= r_data[14693];
                
                r_data[14695] <= r_data[14694];
                
                r_data[14696] <= r_data[14695];
                
                r_data[14697] <= r_data[14696];
                
                r_data[14698] <= r_data[14697];
                
                r_data[14699] <= r_data[14698];
                
                r_data[14700] <= r_data[14699];
                
                r_data[14701] <= r_data[14700];
                
                r_data[14702] <= r_data[14701];
                
                r_data[14703] <= r_data[14702];
                
                r_data[14704] <= r_data[14703];
                
                r_data[14705] <= r_data[14704];
                
                r_data[14706] <= r_data[14705];
                
                r_data[14707] <= r_data[14706];
                
                r_data[14708] <= r_data[14707];
                
                r_data[14709] <= r_data[14708];
                
                r_data[14710] <= r_data[14709];
                
                r_data[14711] <= r_data[14710];
                
                r_data[14712] <= r_data[14711];
                
                r_data[14713] <= r_data[14712];
                
                r_data[14714] <= r_data[14713];
                
                r_data[14715] <= r_data[14714];
                
                r_data[14716] <= r_data[14715];
                
                r_data[14717] <= r_data[14716];
                
                r_data[14718] <= r_data[14717];
                
                r_data[14719] <= r_data[14718];
                
                r_data[14720] <= r_data[14719];
                
                r_data[14721] <= r_data[14720];
                
                r_data[14722] <= r_data[14721];
                
                r_data[14723] <= r_data[14722];
                
                r_data[14724] <= r_data[14723];
                
                r_data[14725] <= r_data[14724];
                
                r_data[14726] <= r_data[14725];
                
                r_data[14727] <= r_data[14726];
                
                r_data[14728] <= r_data[14727];
                
                r_data[14729] <= r_data[14728];
                
                r_data[14730] <= r_data[14729];
                
                r_data[14731] <= r_data[14730];
                
                r_data[14732] <= r_data[14731];
                
                r_data[14733] <= r_data[14732];
                
                r_data[14734] <= r_data[14733];
                
                r_data[14735] <= r_data[14734];
                
                r_data[14736] <= r_data[14735];
                
                r_data[14737] <= r_data[14736];
                
                r_data[14738] <= r_data[14737];
                
                r_data[14739] <= r_data[14738];
                
                r_data[14740] <= r_data[14739];
                
                r_data[14741] <= r_data[14740];
                
                r_data[14742] <= r_data[14741];
                
                r_data[14743] <= r_data[14742];
                
                r_data[14744] <= r_data[14743];
                
                r_data[14745] <= r_data[14744];
                
                r_data[14746] <= r_data[14745];
                
                r_data[14747] <= r_data[14746];
                
                r_data[14748] <= r_data[14747];
                
                r_data[14749] <= r_data[14748];
                
                r_data[14750] <= r_data[14749];
                
                r_data[14751] <= r_data[14750];
                
                r_data[14752] <= r_data[14751];
                
                r_data[14753] <= r_data[14752];
                
                r_data[14754] <= r_data[14753];
                
                r_data[14755] <= r_data[14754];
                
                r_data[14756] <= r_data[14755];
                
                r_data[14757] <= r_data[14756];
                
                r_data[14758] <= r_data[14757];
                
                r_data[14759] <= r_data[14758];
                
                r_data[14760] <= r_data[14759];
                
                r_data[14761] <= r_data[14760];
                
                r_data[14762] <= r_data[14761];
                
                r_data[14763] <= r_data[14762];
                
                r_data[14764] <= r_data[14763];
                
                r_data[14765] <= r_data[14764];
                
                r_data[14766] <= r_data[14765];
                
                r_data[14767] <= r_data[14766];
                
                r_data[14768] <= r_data[14767];
                
                r_data[14769] <= r_data[14768];
                
                r_data[14770] <= r_data[14769];
                
                r_data[14771] <= r_data[14770];
                
                r_data[14772] <= r_data[14771];
                
                r_data[14773] <= r_data[14772];
                
                r_data[14774] <= r_data[14773];
                
                r_data[14775] <= r_data[14774];
                
                r_data[14776] <= r_data[14775];
                
                r_data[14777] <= r_data[14776];
                
                r_data[14778] <= r_data[14777];
                
                r_data[14779] <= r_data[14778];
                
                r_data[14780] <= r_data[14779];
                
                r_data[14781] <= r_data[14780];
                
                r_data[14782] <= r_data[14781];
                
                r_data[14783] <= r_data[14782];
                
                r_data[14784] <= r_data[14783];
                
                r_data[14785] <= r_data[14784];
                
                r_data[14786] <= r_data[14785];
                
                r_data[14787] <= r_data[14786];
                
                r_data[14788] <= r_data[14787];
                
                r_data[14789] <= r_data[14788];
                
                r_data[14790] <= r_data[14789];
                
                r_data[14791] <= r_data[14790];
                
                r_data[14792] <= r_data[14791];
                
                r_data[14793] <= r_data[14792];
                
                r_data[14794] <= r_data[14793];
                
                r_data[14795] <= r_data[14794];
                
                r_data[14796] <= r_data[14795];
                
                r_data[14797] <= r_data[14796];
                
                r_data[14798] <= r_data[14797];
                
                r_data[14799] <= r_data[14798];
                
                r_data[14800] <= r_data[14799];
                
                r_data[14801] <= r_data[14800];
                
                r_data[14802] <= r_data[14801];
                
                r_data[14803] <= r_data[14802];
                
                r_data[14804] <= r_data[14803];
                
                r_data[14805] <= r_data[14804];
                
                r_data[14806] <= r_data[14805];
                
                r_data[14807] <= r_data[14806];
                
                r_data[14808] <= r_data[14807];
                
                r_data[14809] <= r_data[14808];
                
                r_data[14810] <= r_data[14809];
                
                r_data[14811] <= r_data[14810];
                
                r_data[14812] <= r_data[14811];
                
                r_data[14813] <= r_data[14812];
                
                r_data[14814] <= r_data[14813];
                
                r_data[14815] <= r_data[14814];
                
                r_data[14816] <= r_data[14815];
                
                r_data[14817] <= r_data[14816];
                
                r_data[14818] <= r_data[14817];
                
                r_data[14819] <= r_data[14818];
                
                r_data[14820] <= r_data[14819];
                
                r_data[14821] <= r_data[14820];
                
                r_data[14822] <= r_data[14821];
                
                r_data[14823] <= r_data[14822];
                
                r_data[14824] <= r_data[14823];
                
                r_data[14825] <= r_data[14824];
                
                r_data[14826] <= r_data[14825];
                
                r_data[14827] <= r_data[14826];
                
                r_data[14828] <= r_data[14827];
                
                r_data[14829] <= r_data[14828];
                
                r_data[14830] <= r_data[14829];
                
                r_data[14831] <= r_data[14830];
                
                r_data[14832] <= r_data[14831];
                
                r_data[14833] <= r_data[14832];
                
                r_data[14834] <= r_data[14833];
                
                r_data[14835] <= r_data[14834];
                
                r_data[14836] <= r_data[14835];
                
                r_data[14837] <= r_data[14836];
                
                r_data[14838] <= r_data[14837];
                
                r_data[14839] <= r_data[14838];
                
                r_data[14840] <= r_data[14839];
                
                r_data[14841] <= r_data[14840];
                
                r_data[14842] <= r_data[14841];
                
                r_data[14843] <= r_data[14842];
                
                r_data[14844] <= r_data[14843];
                
                r_data[14845] <= r_data[14844];
                
                r_data[14846] <= r_data[14845];
                
                r_data[14847] <= r_data[14846];
                
                r_data[14848] <= r_data[14847];
                
                r_data[14849] <= r_data[14848];
                
                r_data[14850] <= r_data[14849];
                
                r_data[14851] <= r_data[14850];
                
                r_data[14852] <= r_data[14851];
                
                r_data[14853] <= r_data[14852];
                
                r_data[14854] <= r_data[14853];
                
                r_data[14855] <= r_data[14854];
                
                r_data[14856] <= r_data[14855];
                
                r_data[14857] <= r_data[14856];
                
                r_data[14858] <= r_data[14857];
                
                r_data[14859] <= r_data[14858];
                
                r_data[14860] <= r_data[14859];
                
                r_data[14861] <= r_data[14860];
                
                r_data[14862] <= r_data[14861];
                
                r_data[14863] <= r_data[14862];
                
                r_data[14864] <= r_data[14863];
                
                r_data[14865] <= r_data[14864];
                
                r_data[14866] <= r_data[14865];
                
                r_data[14867] <= r_data[14866];
                
                r_data[14868] <= r_data[14867];
                
                r_data[14869] <= r_data[14868];
                
                r_data[14870] <= r_data[14869];
                
                r_data[14871] <= r_data[14870];
                
                r_data[14872] <= r_data[14871];
                
                r_data[14873] <= r_data[14872];
                
                r_data[14874] <= r_data[14873];
                
                r_data[14875] <= r_data[14874];
                
                r_data[14876] <= r_data[14875];
                
                r_data[14877] <= r_data[14876];
                
                r_data[14878] <= r_data[14877];
                
                r_data[14879] <= r_data[14878];
                
                r_data[14880] <= r_data[14879];
                
                r_data[14881] <= r_data[14880];
                
                r_data[14882] <= r_data[14881];
                
                r_data[14883] <= r_data[14882];
                
                r_data[14884] <= r_data[14883];
                
                r_data[14885] <= r_data[14884];
                
                r_data[14886] <= r_data[14885];
                
                r_data[14887] <= r_data[14886];
                
                r_data[14888] <= r_data[14887];
                
                r_data[14889] <= r_data[14888];
                
                r_data[14890] <= r_data[14889];
                
                r_data[14891] <= r_data[14890];
                
                r_data[14892] <= r_data[14891];
                
                r_data[14893] <= r_data[14892];
                
                r_data[14894] <= r_data[14893];
                
                r_data[14895] <= r_data[14894];
                
                r_data[14896] <= r_data[14895];
                
                r_data[14897] <= r_data[14896];
                
                r_data[14898] <= r_data[14897];
                
                r_data[14899] <= r_data[14898];
                
                r_data[14900] <= r_data[14899];
                
                r_data[14901] <= r_data[14900];
                
                r_data[14902] <= r_data[14901];
                
                r_data[14903] <= r_data[14902];
                
                r_data[14904] <= r_data[14903];
                
                r_data[14905] <= r_data[14904];
                
                r_data[14906] <= r_data[14905];
                
                r_data[14907] <= r_data[14906];
                
                r_data[14908] <= r_data[14907];
                
                r_data[14909] <= r_data[14908];
                
                r_data[14910] <= r_data[14909];
                
                r_data[14911] <= r_data[14910];
                
                r_data[14912] <= r_data[14911];
                
                r_data[14913] <= r_data[14912];
                
                r_data[14914] <= r_data[14913];
                
                r_data[14915] <= r_data[14914];
                
                r_data[14916] <= r_data[14915];
                
                r_data[14917] <= r_data[14916];
                
                r_data[14918] <= r_data[14917];
                
                r_data[14919] <= r_data[14918];
                
                r_data[14920] <= r_data[14919];
                
                r_data[14921] <= r_data[14920];
                
                r_data[14922] <= r_data[14921];
                
                r_data[14923] <= r_data[14922];
                
                r_data[14924] <= r_data[14923];
                
                r_data[14925] <= r_data[14924];
                
                r_data[14926] <= r_data[14925];
                
                r_data[14927] <= r_data[14926];
                
                r_data[14928] <= r_data[14927];
                
                r_data[14929] <= r_data[14928];
                
                r_data[14930] <= r_data[14929];
                
                r_data[14931] <= r_data[14930];
                
                r_data[14932] <= r_data[14931];
                
                r_data[14933] <= r_data[14932];
                
                r_data[14934] <= r_data[14933];
                
                r_data[14935] <= r_data[14934];
                
                r_data[14936] <= r_data[14935];
                
                r_data[14937] <= r_data[14936];
                
                r_data[14938] <= r_data[14937];
                
                r_data[14939] <= r_data[14938];
                
                r_data[14940] <= r_data[14939];
                
                r_data[14941] <= r_data[14940];
                
                r_data[14942] <= r_data[14941];
                
                r_data[14943] <= r_data[14942];
                
                r_data[14944] <= r_data[14943];
                
                r_data[14945] <= r_data[14944];
                
                r_data[14946] <= r_data[14945];
                
                r_data[14947] <= r_data[14946];
                
                r_data[14948] <= r_data[14947];
                
                r_data[14949] <= r_data[14948];
                
                r_data[14950] <= r_data[14949];
                
                r_data[14951] <= r_data[14950];
                
                r_data[14952] <= r_data[14951];
                
                r_data[14953] <= r_data[14952];
                
                r_data[14954] <= r_data[14953];
                
                r_data[14955] <= r_data[14954];
                
                r_data[14956] <= r_data[14955];
                
                r_data[14957] <= r_data[14956];
                
                r_data[14958] <= r_data[14957];
                
                r_data[14959] <= r_data[14958];
                
                r_data[14960] <= r_data[14959];
                
                r_data[14961] <= r_data[14960];
                
                r_data[14962] <= r_data[14961];
                
                r_data[14963] <= r_data[14962];
                
                r_data[14964] <= r_data[14963];
                
                r_data[14965] <= r_data[14964];
                
                r_data[14966] <= r_data[14965];
                
                r_data[14967] <= r_data[14966];
                
                r_data[14968] <= r_data[14967];
                
                r_data[14969] <= r_data[14968];
                
                r_data[14970] <= r_data[14969];
                
                r_data[14971] <= r_data[14970];
                
                r_data[14972] <= r_data[14971];
                
                r_data[14973] <= r_data[14972];
                
                r_data[14974] <= r_data[14973];
                
                r_data[14975] <= r_data[14974];
                
                r_data[14976] <= r_data[14975];
                
                r_data[14977] <= r_data[14976];
                
                r_data[14978] <= r_data[14977];
                
                r_data[14979] <= r_data[14978];
                
                r_data[14980] <= r_data[14979];
                
                r_data[14981] <= r_data[14980];
                
                r_data[14982] <= r_data[14981];
                
                r_data[14983] <= r_data[14982];
                
                r_data[14984] <= r_data[14983];
                
                r_data[14985] <= r_data[14984];
                
                r_data[14986] <= r_data[14985];
                
                r_data[14987] <= r_data[14986];
                
                r_data[14988] <= r_data[14987];
                
                r_data[14989] <= r_data[14988];
                
                r_data[14990] <= r_data[14989];
                
                r_data[14991] <= r_data[14990];
                
                r_data[14992] <= r_data[14991];
                
                r_data[14993] <= r_data[14992];
                
                r_data[14994] <= r_data[14993];
                
                r_data[14995] <= r_data[14994];
                
                r_data[14996] <= r_data[14995];
                
                r_data[14997] <= r_data[14996];
                
                r_data[14998] <= r_data[14997];
                
                r_data[14999] <= r_data[14998];
                
                r_data[15000] <= r_data[14999];
                
                r_data[15001] <= r_data[15000];
                
                r_data[15002] <= r_data[15001];
                
                r_data[15003] <= r_data[15002];
                
                r_data[15004] <= r_data[15003];
                
                r_data[15005] <= r_data[15004];
                
                r_data[15006] <= r_data[15005];
                
                r_data[15007] <= r_data[15006];
                
                r_data[15008] <= r_data[15007];
                
                r_data[15009] <= r_data[15008];
                
                r_data[15010] <= r_data[15009];
                
                r_data[15011] <= r_data[15010];
                
                r_data[15012] <= r_data[15011];
                
                r_data[15013] <= r_data[15012];
                
                r_data[15014] <= r_data[15013];
                
                r_data[15015] <= r_data[15014];
                
                r_data[15016] <= r_data[15015];
                
                r_data[15017] <= r_data[15016];
                
                r_data[15018] <= r_data[15017];
                
                r_data[15019] <= r_data[15018];
                
                r_data[15020] <= r_data[15019];
                
                r_data[15021] <= r_data[15020];
                
                r_data[15022] <= r_data[15021];
                
                r_data[15023] <= r_data[15022];
                
                r_data[15024] <= r_data[15023];
                
                r_data[15025] <= r_data[15024];
                
                r_data[15026] <= r_data[15025];
                
                r_data[15027] <= r_data[15026];
                
                r_data[15028] <= r_data[15027];
                
                r_data[15029] <= r_data[15028];
                
                r_data[15030] <= r_data[15029];
                
                r_data[15031] <= r_data[15030];
                
                r_data[15032] <= r_data[15031];
                
                r_data[15033] <= r_data[15032];
                
                r_data[15034] <= r_data[15033];
                
                r_data[15035] <= r_data[15034];
                
                r_data[15036] <= r_data[15035];
                
                r_data[15037] <= r_data[15036];
                
                r_data[15038] <= r_data[15037];
                
                r_data[15039] <= r_data[15038];
                
                r_data[15040] <= r_data[15039];
                
                r_data[15041] <= r_data[15040];
                
                r_data[15042] <= r_data[15041];
                
                r_data[15043] <= r_data[15042];
                
                r_data[15044] <= r_data[15043];
                
                r_data[15045] <= r_data[15044];
                
                r_data[15046] <= r_data[15045];
                
                r_data[15047] <= r_data[15046];
                
                r_data[15048] <= r_data[15047];
                
                r_data[15049] <= r_data[15048];
                
                r_data[15050] <= r_data[15049];
                
                r_data[15051] <= r_data[15050];
                
                r_data[15052] <= r_data[15051];
                
                r_data[15053] <= r_data[15052];
                
                r_data[15054] <= r_data[15053];
                
                r_data[15055] <= r_data[15054];
                
                r_data[15056] <= r_data[15055];
                
                r_data[15057] <= r_data[15056];
                
                r_data[15058] <= r_data[15057];
                
                r_data[15059] <= r_data[15058];
                
                r_data[15060] <= r_data[15059];
                
                r_data[15061] <= r_data[15060];
                
                r_data[15062] <= r_data[15061];
                
                r_data[15063] <= r_data[15062];
                
                r_data[15064] <= r_data[15063];
                
                r_data[15065] <= r_data[15064];
                
                r_data[15066] <= r_data[15065];
                
                r_data[15067] <= r_data[15066];
                
                r_data[15068] <= r_data[15067];
                
                r_data[15069] <= r_data[15068];
                
                r_data[15070] <= r_data[15069];
                
                r_data[15071] <= r_data[15070];
                
                r_data[15072] <= r_data[15071];
                
                r_data[15073] <= r_data[15072];
                
                r_data[15074] <= r_data[15073];
                
                r_data[15075] <= r_data[15074];
                
                r_data[15076] <= r_data[15075];
                
                r_data[15077] <= r_data[15076];
                
                r_data[15078] <= r_data[15077];
                
                r_data[15079] <= r_data[15078];
                
                r_data[15080] <= r_data[15079];
                
                r_data[15081] <= r_data[15080];
                
                r_data[15082] <= r_data[15081];
                
                r_data[15083] <= r_data[15082];
                
                r_data[15084] <= r_data[15083];
                
                r_data[15085] <= r_data[15084];
                
                r_data[15086] <= r_data[15085];
                
                r_data[15087] <= r_data[15086];
                
                r_data[15088] <= r_data[15087];
                
                r_data[15089] <= r_data[15088];
                
                r_data[15090] <= r_data[15089];
                
                r_data[15091] <= r_data[15090];
                
                r_data[15092] <= r_data[15091];
                
                r_data[15093] <= r_data[15092];
                
                r_data[15094] <= r_data[15093];
                
                r_data[15095] <= r_data[15094];
                
                r_data[15096] <= r_data[15095];
                
                r_data[15097] <= r_data[15096];
                
                r_data[15098] <= r_data[15097];
                
                r_data[15099] <= r_data[15098];
                
                r_data[15100] <= r_data[15099];
                
                r_data[15101] <= r_data[15100];
                
                r_data[15102] <= r_data[15101];
                
                r_data[15103] <= r_data[15102];
                
                r_data[15104] <= r_data[15103];
                
                r_data[15105] <= r_data[15104];
                
                r_data[15106] <= r_data[15105];
                
                r_data[15107] <= r_data[15106];
                
                r_data[15108] <= r_data[15107];
                
                r_data[15109] <= r_data[15108];
                
                r_data[15110] <= r_data[15109];
                
                r_data[15111] <= r_data[15110];
                
                r_data[15112] <= r_data[15111];
                
                r_data[15113] <= r_data[15112];
                
                r_data[15114] <= r_data[15113];
                
                r_data[15115] <= r_data[15114];
                
                r_data[15116] <= r_data[15115];
                
                r_data[15117] <= r_data[15116];
                
                r_data[15118] <= r_data[15117];
                
                r_data[15119] <= r_data[15118];
                
                r_data[15120] <= r_data[15119];
                
                r_data[15121] <= r_data[15120];
                
                r_data[15122] <= r_data[15121];
                
                r_data[15123] <= r_data[15122];
                
                r_data[15124] <= r_data[15123];
                
                r_data[15125] <= r_data[15124];
                
                r_data[15126] <= r_data[15125];
                
                r_data[15127] <= r_data[15126];
                
                r_data[15128] <= r_data[15127];
                
                r_data[15129] <= r_data[15128];
                
                r_data[15130] <= r_data[15129];
                
                r_data[15131] <= r_data[15130];
                
                r_data[15132] <= r_data[15131];
                
                r_data[15133] <= r_data[15132];
                
                r_data[15134] <= r_data[15133];
                
                r_data[15135] <= r_data[15134];
                
                r_data[15136] <= r_data[15135];
                
                r_data[15137] <= r_data[15136];
                
                r_data[15138] <= r_data[15137];
                
                r_data[15139] <= r_data[15138];
                
                r_data[15140] <= r_data[15139];
                
                r_data[15141] <= r_data[15140];
                
                r_data[15142] <= r_data[15141];
                
                r_data[15143] <= r_data[15142];
                
                r_data[15144] <= r_data[15143];
                
                r_data[15145] <= r_data[15144];
                
                r_data[15146] <= r_data[15145];
                
                r_data[15147] <= r_data[15146];
                
                r_data[15148] <= r_data[15147];
                
                r_data[15149] <= r_data[15148];
                
                r_data[15150] <= r_data[15149];
                
                r_data[15151] <= r_data[15150];
                
                r_data[15152] <= r_data[15151];
                
                r_data[15153] <= r_data[15152];
                
                r_data[15154] <= r_data[15153];
                
                r_data[15155] <= r_data[15154];
                
                r_data[15156] <= r_data[15155];
                
                r_data[15157] <= r_data[15156];
                
                r_data[15158] <= r_data[15157];
                
                r_data[15159] <= r_data[15158];
                
                r_data[15160] <= r_data[15159];
                
                r_data[15161] <= r_data[15160];
                
                r_data[15162] <= r_data[15161];
                
                r_data[15163] <= r_data[15162];
                
                r_data[15164] <= r_data[15163];
                
                r_data[15165] <= r_data[15164];
                
                r_data[15166] <= r_data[15165];
                
                r_data[15167] <= r_data[15166];
                
                r_data[15168] <= r_data[15167];
                
                r_data[15169] <= r_data[15168];
                
                r_data[15170] <= r_data[15169];
                
                r_data[15171] <= r_data[15170];
                
                r_data[15172] <= r_data[15171];
                
                r_data[15173] <= r_data[15172];
                
                r_data[15174] <= r_data[15173];
                
                r_data[15175] <= r_data[15174];
                
                r_data[15176] <= r_data[15175];
                
                r_data[15177] <= r_data[15176];
                
                r_data[15178] <= r_data[15177];
                
                r_data[15179] <= r_data[15178];
                
                r_data[15180] <= r_data[15179];
                
                r_data[15181] <= r_data[15180];
                
                r_data[15182] <= r_data[15181];
                
                r_data[15183] <= r_data[15182];
                
                r_data[15184] <= r_data[15183];
                
                r_data[15185] <= r_data[15184];
                
                r_data[15186] <= r_data[15185];
                
                r_data[15187] <= r_data[15186];
                
                r_data[15188] <= r_data[15187];
                
                r_data[15189] <= r_data[15188];
                
                r_data[15190] <= r_data[15189];
                
                r_data[15191] <= r_data[15190];
                
                r_data[15192] <= r_data[15191];
                
                r_data[15193] <= r_data[15192];
                
                r_data[15194] <= r_data[15193];
                
                r_data[15195] <= r_data[15194];
                
                r_data[15196] <= r_data[15195];
                
                r_data[15197] <= r_data[15196];
                
                r_data[15198] <= r_data[15197];
                
                r_data[15199] <= r_data[15198];
                
                r_data[15200] <= r_data[15199];
                
                r_data[15201] <= r_data[15200];
                
                r_data[15202] <= r_data[15201];
                
                r_data[15203] <= r_data[15202];
                
                r_data[15204] <= r_data[15203];
                
                r_data[15205] <= r_data[15204];
                
                r_data[15206] <= r_data[15205];
                
                r_data[15207] <= r_data[15206];
                
                r_data[15208] <= r_data[15207];
                
                r_data[15209] <= r_data[15208];
                
                r_data[15210] <= r_data[15209];
                
                r_data[15211] <= r_data[15210];
                
                r_data[15212] <= r_data[15211];
                
                r_data[15213] <= r_data[15212];
                
                r_data[15214] <= r_data[15213];
                
                r_data[15215] <= r_data[15214];
                
                r_data[15216] <= r_data[15215];
                
                r_data[15217] <= r_data[15216];
                
                r_data[15218] <= r_data[15217];
                
                r_data[15219] <= r_data[15218];
                
                r_data[15220] <= r_data[15219];
                
                r_data[15221] <= r_data[15220];
                
                r_data[15222] <= r_data[15221];
                
                r_data[15223] <= r_data[15222];
                
                r_data[15224] <= r_data[15223];
                
                r_data[15225] <= r_data[15224];
                
                r_data[15226] <= r_data[15225];
                
                r_data[15227] <= r_data[15226];
                
                r_data[15228] <= r_data[15227];
                
                r_data[15229] <= r_data[15228];
                
                r_data[15230] <= r_data[15229];
                
                r_data[15231] <= r_data[15230];
                
                r_data[15232] <= r_data[15231];
                
                r_data[15233] <= r_data[15232];
                
                r_data[15234] <= r_data[15233];
                
                r_data[15235] <= r_data[15234];
                
                r_data[15236] <= r_data[15235];
                
                r_data[15237] <= r_data[15236];
                
                r_data[15238] <= r_data[15237];
                
                r_data[15239] <= r_data[15238];
                
                r_data[15240] <= r_data[15239];
                
                r_data[15241] <= r_data[15240];
                
                r_data[15242] <= r_data[15241];
                
                r_data[15243] <= r_data[15242];
                
                r_data[15244] <= r_data[15243];
                
                r_data[15245] <= r_data[15244];
                
                r_data[15246] <= r_data[15245];
                
                r_data[15247] <= r_data[15246];
                
                r_data[15248] <= r_data[15247];
                
                r_data[15249] <= r_data[15248];
                
                r_data[15250] <= r_data[15249];
                
                r_data[15251] <= r_data[15250];
                
                r_data[15252] <= r_data[15251];
                
                r_data[15253] <= r_data[15252];
                
                r_data[15254] <= r_data[15253];
                
                r_data[15255] <= r_data[15254];
                
                r_data[15256] <= r_data[15255];
                
                r_data[15257] <= r_data[15256];
                
                r_data[15258] <= r_data[15257];
                
                r_data[15259] <= r_data[15258];
                
                r_data[15260] <= r_data[15259];
                
                r_data[15261] <= r_data[15260];
                
                r_data[15262] <= r_data[15261];
                
                r_data[15263] <= r_data[15262];
                
                r_data[15264] <= r_data[15263];
                
                r_data[15265] <= r_data[15264];
                
                r_data[15266] <= r_data[15265];
                
                r_data[15267] <= r_data[15266];
                
                r_data[15268] <= r_data[15267];
                
                r_data[15269] <= r_data[15268];
                
                r_data[15270] <= r_data[15269];
                
                r_data[15271] <= r_data[15270];
                
                r_data[15272] <= r_data[15271];
                
                r_data[15273] <= r_data[15272];
                
                r_data[15274] <= r_data[15273];
                
                r_data[15275] <= r_data[15274];
                
                r_data[15276] <= r_data[15275];
                
                r_data[15277] <= r_data[15276];
                
                r_data[15278] <= r_data[15277];
                
                r_data[15279] <= r_data[15278];
                
                r_data[15280] <= r_data[15279];
                
                r_data[15281] <= r_data[15280];
                
                r_data[15282] <= r_data[15281];
                
                r_data[15283] <= r_data[15282];
                
                r_data[15284] <= r_data[15283];
                
                r_data[15285] <= r_data[15284];
                
                r_data[15286] <= r_data[15285];
                
                r_data[15287] <= r_data[15286];
                
                r_data[15288] <= r_data[15287];
                
                r_data[15289] <= r_data[15288];
                
                r_data[15290] <= r_data[15289];
                
                r_data[15291] <= r_data[15290];
                
                r_data[15292] <= r_data[15291];
                
                r_data[15293] <= r_data[15292];
                
                r_data[15294] <= r_data[15293];
                
                r_data[15295] <= r_data[15294];
                
                r_data[15296] <= r_data[15295];
                
                r_data[15297] <= r_data[15296];
                
                r_data[15298] <= r_data[15297];
                
                r_data[15299] <= r_data[15298];
                
                r_data[15300] <= r_data[15299];
                
                r_data[15301] <= r_data[15300];
                
                r_data[15302] <= r_data[15301];
                
                r_data[15303] <= r_data[15302];
                
                r_data[15304] <= r_data[15303];
                
                r_data[15305] <= r_data[15304];
                
                r_data[15306] <= r_data[15305];
                
                r_data[15307] <= r_data[15306];
                
                r_data[15308] <= r_data[15307];
                
                r_data[15309] <= r_data[15308];
                
                r_data[15310] <= r_data[15309];
                
                r_data[15311] <= r_data[15310];
                
                r_data[15312] <= r_data[15311];
                
                r_data[15313] <= r_data[15312];
                
                r_data[15314] <= r_data[15313];
                
                r_data[15315] <= r_data[15314];
                
                r_data[15316] <= r_data[15315];
                
                r_data[15317] <= r_data[15316];
                
                r_data[15318] <= r_data[15317];
                
                r_data[15319] <= r_data[15318];
                
                r_data[15320] <= r_data[15319];
                
                r_data[15321] <= r_data[15320];
                
                r_data[15322] <= r_data[15321];
                
                r_data[15323] <= r_data[15322];
                
                r_data[15324] <= r_data[15323];
                
                r_data[15325] <= r_data[15324];
                
                r_data[15326] <= r_data[15325];
                
                r_data[15327] <= r_data[15326];
                
                r_data[15328] <= r_data[15327];
                
                r_data[15329] <= r_data[15328];
                
                r_data[15330] <= r_data[15329];
                
                r_data[15331] <= r_data[15330];
                
                r_data[15332] <= r_data[15331];
                
                r_data[15333] <= r_data[15332];
                
                r_data[15334] <= r_data[15333];
                
                r_data[15335] <= r_data[15334];
                
                r_data[15336] <= r_data[15335];
                
                r_data[15337] <= r_data[15336];
                
                r_data[15338] <= r_data[15337];
                
                r_data[15339] <= r_data[15338];
                
                r_data[15340] <= r_data[15339];
                
                r_data[15341] <= r_data[15340];
                
                r_data[15342] <= r_data[15341];
                
                r_data[15343] <= r_data[15342];
                
                r_data[15344] <= r_data[15343];
                
                r_data[15345] <= r_data[15344];
                
                r_data[15346] <= r_data[15345];
                
                r_data[15347] <= r_data[15346];
                
                r_data[15348] <= r_data[15347];
                
                r_data[15349] <= r_data[15348];
                
                r_data[15350] <= r_data[15349];
                
                r_data[15351] <= r_data[15350];
                
                r_data[15352] <= r_data[15351];
                
                r_data[15353] <= r_data[15352];
                
                r_data[15354] <= r_data[15353];
                
                r_data[15355] <= r_data[15354];
                
                r_data[15356] <= r_data[15355];
                
                r_data[15357] <= r_data[15356];
                
                r_data[15358] <= r_data[15357];
                
                r_data[15359] <= r_data[15358];
                
                r_data[15360] <= r_data[15359];
                
                r_data[15361] <= r_data[15360];
                
                r_data[15362] <= r_data[15361];
                
                r_data[15363] <= r_data[15362];
                
                r_data[15364] <= r_data[15363];
                
                r_data[15365] <= r_data[15364];
                
                r_data[15366] <= r_data[15365];
                
                r_data[15367] <= r_data[15366];
                
                r_data[15368] <= r_data[15367];
                
                r_data[15369] <= r_data[15368];
                
                r_data[15370] <= r_data[15369];
                
                r_data[15371] <= r_data[15370];
                
                r_data[15372] <= r_data[15371];
                
                r_data[15373] <= r_data[15372];
                
                r_data[15374] <= r_data[15373];
                
                r_data[15375] <= r_data[15374];
                
                r_data[15376] <= r_data[15375];
                
                r_data[15377] <= r_data[15376];
                
                r_data[15378] <= r_data[15377];
                
                r_data[15379] <= r_data[15378];
                
                r_data[15380] <= r_data[15379];
                
                r_data[15381] <= r_data[15380];
                
                r_data[15382] <= r_data[15381];
                
                r_data[15383] <= r_data[15382];
                
                r_data[15384] <= r_data[15383];
                
                r_data[15385] <= r_data[15384];
                
                r_data[15386] <= r_data[15385];
                
                r_data[15387] <= r_data[15386];
                
                r_data[15388] <= r_data[15387];
                
                r_data[15389] <= r_data[15388];
                
                r_data[15390] <= r_data[15389];
                
                r_data[15391] <= r_data[15390];
                
                r_data[15392] <= r_data[15391];
                
                r_data[15393] <= r_data[15392];
                
                r_data[15394] <= r_data[15393];
                
                r_data[15395] <= r_data[15394];
                
                r_data[15396] <= r_data[15395];
                
                r_data[15397] <= r_data[15396];
                
                r_data[15398] <= r_data[15397];
                
                r_data[15399] <= r_data[15398];
                
                r_data[15400] <= r_data[15399];
                
                r_data[15401] <= r_data[15400];
                
                r_data[15402] <= r_data[15401];
                
                r_data[15403] <= r_data[15402];
                
                r_data[15404] <= r_data[15403];
                
                r_data[15405] <= r_data[15404];
                
                r_data[15406] <= r_data[15405];
                
                r_data[15407] <= r_data[15406];
                
                r_data[15408] <= r_data[15407];
                
                r_data[15409] <= r_data[15408];
                
                r_data[15410] <= r_data[15409];
                
                r_data[15411] <= r_data[15410];
                
                r_data[15412] <= r_data[15411];
                
                r_data[15413] <= r_data[15412];
                
                r_data[15414] <= r_data[15413];
                
                r_data[15415] <= r_data[15414];
                
                r_data[15416] <= r_data[15415];
                
                r_data[15417] <= r_data[15416];
                
                r_data[15418] <= r_data[15417];
                
                r_data[15419] <= r_data[15418];
                
                r_data[15420] <= r_data[15419];
                
                r_data[15421] <= r_data[15420];
                
                r_data[15422] <= r_data[15421];
                
                r_data[15423] <= r_data[15422];
                
                r_data[15424] <= r_data[15423];
                
                r_data[15425] <= r_data[15424];
                
                r_data[15426] <= r_data[15425];
                
                r_data[15427] <= r_data[15426];
                
                r_data[15428] <= r_data[15427];
                
                r_data[15429] <= r_data[15428];
                
                r_data[15430] <= r_data[15429];
                
                r_data[15431] <= r_data[15430];
                
                r_data[15432] <= r_data[15431];
                
                r_data[15433] <= r_data[15432];
                
                r_data[15434] <= r_data[15433];
                
                r_data[15435] <= r_data[15434];
                
                r_data[15436] <= r_data[15435];
                
                r_data[15437] <= r_data[15436];
                
                r_data[15438] <= r_data[15437];
                
                r_data[15439] <= r_data[15438];
                
                r_data[15440] <= r_data[15439];
                
                r_data[15441] <= r_data[15440];
                
                r_data[15442] <= r_data[15441];
                
                r_data[15443] <= r_data[15442];
                
                r_data[15444] <= r_data[15443];
                
                r_data[15445] <= r_data[15444];
                
                r_data[15446] <= r_data[15445];
                
                r_data[15447] <= r_data[15446];
                
                r_data[15448] <= r_data[15447];
                
                r_data[15449] <= r_data[15448];
                
                r_data[15450] <= r_data[15449];
                
                r_data[15451] <= r_data[15450];
                
                r_data[15452] <= r_data[15451];
                
                r_data[15453] <= r_data[15452];
                
                r_data[15454] <= r_data[15453];
                
                r_data[15455] <= r_data[15454];
                
                r_data[15456] <= r_data[15455];
                
                r_data[15457] <= r_data[15456];
                
                r_data[15458] <= r_data[15457];
                
                r_data[15459] <= r_data[15458];
                
                r_data[15460] <= r_data[15459];
                
                r_data[15461] <= r_data[15460];
                
                r_data[15462] <= r_data[15461];
                
                r_data[15463] <= r_data[15462];
                
                r_data[15464] <= r_data[15463];
                
                r_data[15465] <= r_data[15464];
                
                r_data[15466] <= r_data[15465];
                
                r_data[15467] <= r_data[15466];
                
                r_data[15468] <= r_data[15467];
                
                r_data[15469] <= r_data[15468];
                
                r_data[15470] <= r_data[15469];
                
                r_data[15471] <= r_data[15470];
                
                r_data[15472] <= r_data[15471];
                
                r_data[15473] <= r_data[15472];
                
                r_data[15474] <= r_data[15473];
                
                r_data[15475] <= r_data[15474];
                
                r_data[15476] <= r_data[15475];
                
                r_data[15477] <= r_data[15476];
                
                r_data[15478] <= r_data[15477];
                
                r_data[15479] <= r_data[15478];
                
                r_data[15480] <= r_data[15479];
                
                r_data[15481] <= r_data[15480];
                
                r_data[15482] <= r_data[15481];
                
                r_data[15483] <= r_data[15482];
                
                r_data[15484] <= r_data[15483];
                
                r_data[15485] <= r_data[15484];
                
                r_data[15486] <= r_data[15485];
                
                r_data[15487] <= r_data[15486];
                
                r_data[15488] <= r_data[15487];
                
                r_data[15489] <= r_data[15488];
                
                r_data[15490] <= r_data[15489];
                
                r_data[15491] <= r_data[15490];
                
                r_data[15492] <= r_data[15491];
                
                r_data[15493] <= r_data[15492];
                
                r_data[15494] <= r_data[15493];
                
                r_data[15495] <= r_data[15494];
                
                r_data[15496] <= r_data[15495];
                
                r_data[15497] <= r_data[15496];
                
                r_data[15498] <= r_data[15497];
                
                r_data[15499] <= r_data[15498];
                
                r_data[15500] <= r_data[15499];
                
                r_data[15501] <= r_data[15500];
                
                r_data[15502] <= r_data[15501];
                
                r_data[15503] <= r_data[15502];
                
                r_data[15504] <= r_data[15503];
                
                r_data[15505] <= r_data[15504];
                
                r_data[15506] <= r_data[15505];
                
                r_data[15507] <= r_data[15506];
                
                r_data[15508] <= r_data[15507];
                
                r_data[15509] <= r_data[15508];
                
                r_data[15510] <= r_data[15509];
                
                r_data[15511] <= r_data[15510];
                
                r_data[15512] <= r_data[15511];
                
                r_data[15513] <= r_data[15512];
                
                r_data[15514] <= r_data[15513];
                
                r_data[15515] <= r_data[15514];
                
                r_data[15516] <= r_data[15515];
                
                r_data[15517] <= r_data[15516];
                
                r_data[15518] <= r_data[15517];
                
                r_data[15519] <= r_data[15518];
                
                r_data[15520] <= r_data[15519];
                
                r_data[15521] <= r_data[15520];
                
                r_data[15522] <= r_data[15521];
                
                r_data[15523] <= r_data[15522];
                
                r_data[15524] <= r_data[15523];
                
                r_data[15525] <= r_data[15524];
                
                r_data[15526] <= r_data[15525];
                
                r_data[15527] <= r_data[15526];
                
                r_data[15528] <= r_data[15527];
                
                r_data[15529] <= r_data[15528];
                
                r_data[15530] <= r_data[15529];
                
                r_data[15531] <= r_data[15530];
                
                r_data[15532] <= r_data[15531];
                
                r_data[15533] <= r_data[15532];
                
                r_data[15534] <= r_data[15533];
                
                r_data[15535] <= r_data[15534];
                
                r_data[15536] <= r_data[15535];
                
                r_data[15537] <= r_data[15536];
                
                r_data[15538] <= r_data[15537];
                
                r_data[15539] <= r_data[15538];
                
                r_data[15540] <= r_data[15539];
                
                r_data[15541] <= r_data[15540];
                
                r_data[15542] <= r_data[15541];
                
                r_data[15543] <= r_data[15542];
                
                r_data[15544] <= r_data[15543];
                
                r_data[15545] <= r_data[15544];
                
                r_data[15546] <= r_data[15545];
                
                r_data[15547] <= r_data[15546];
                
                r_data[15548] <= r_data[15547];
                
                r_data[15549] <= r_data[15548];
                
                r_data[15550] <= r_data[15549];
                
                r_data[15551] <= r_data[15550];
                
                r_data[15552] <= r_data[15551];
                
                r_data[15553] <= r_data[15552];
                
                r_data[15554] <= r_data[15553];
                
                r_data[15555] <= r_data[15554];
                
                r_data[15556] <= r_data[15555];
                
                r_data[15557] <= r_data[15556];
                
                r_data[15558] <= r_data[15557];
                
                r_data[15559] <= r_data[15558];
                
                r_data[15560] <= r_data[15559];
                
                r_data[15561] <= r_data[15560];
                
                r_data[15562] <= r_data[15561];
                
                r_data[15563] <= r_data[15562];
                
                r_data[15564] <= r_data[15563];
                
                r_data[15565] <= r_data[15564];
                
                r_data[15566] <= r_data[15565];
                
                r_data[15567] <= r_data[15566];
                
                r_data[15568] <= r_data[15567];
                
                r_data[15569] <= r_data[15568];
                
                r_data[15570] <= r_data[15569];
                
                r_data[15571] <= r_data[15570];
                
                r_data[15572] <= r_data[15571];
                
                r_data[15573] <= r_data[15572];
                
                r_data[15574] <= r_data[15573];
                
                r_data[15575] <= r_data[15574];
                
                r_data[15576] <= r_data[15575];
                
                r_data[15577] <= r_data[15576];
                
                r_data[15578] <= r_data[15577];
                
                r_data[15579] <= r_data[15578];
                
                r_data[15580] <= r_data[15579];
                
                r_data[15581] <= r_data[15580];
                
                r_data[15582] <= r_data[15581];
                
                r_data[15583] <= r_data[15582];
                
                r_data[15584] <= r_data[15583];
                
                r_data[15585] <= r_data[15584];
                
                r_data[15586] <= r_data[15585];
                
                r_data[15587] <= r_data[15586];
                
                r_data[15588] <= r_data[15587];
                
                r_data[15589] <= r_data[15588];
                
                r_data[15590] <= r_data[15589];
                
                r_data[15591] <= r_data[15590];
                
                r_data[15592] <= r_data[15591];
                
                r_data[15593] <= r_data[15592];
                
                r_data[15594] <= r_data[15593];
                
                r_data[15595] <= r_data[15594];
                
                r_data[15596] <= r_data[15595];
                
                r_data[15597] <= r_data[15596];
                
                r_data[15598] <= r_data[15597];
                
                r_data[15599] <= r_data[15598];
                
                r_data[15600] <= r_data[15599];
                
                r_data[15601] <= r_data[15600];
                
                r_data[15602] <= r_data[15601];
                
                r_data[15603] <= r_data[15602];
                
                r_data[15604] <= r_data[15603];
                
                r_data[15605] <= r_data[15604];
                
                r_data[15606] <= r_data[15605];
                
                r_data[15607] <= r_data[15606];
                
                r_data[15608] <= r_data[15607];
                
                r_data[15609] <= r_data[15608];
                
                r_data[15610] <= r_data[15609];
                
                r_data[15611] <= r_data[15610];
                
                r_data[15612] <= r_data[15611];
                
                r_data[15613] <= r_data[15612];
                
                r_data[15614] <= r_data[15613];
                
                r_data[15615] <= r_data[15614];
                
                r_data[15616] <= r_data[15615];
                
                r_data[15617] <= r_data[15616];
                
                r_data[15618] <= r_data[15617];
                
                r_data[15619] <= r_data[15618];
                
                r_data[15620] <= r_data[15619];
                
                r_data[15621] <= r_data[15620];
                
                r_data[15622] <= r_data[15621];
                
                r_data[15623] <= r_data[15622];
                
                r_data[15624] <= r_data[15623];
                
                r_data[15625] <= r_data[15624];
                
                r_data[15626] <= r_data[15625];
                
                r_data[15627] <= r_data[15626];
                
                r_data[15628] <= r_data[15627];
                
                r_data[15629] <= r_data[15628];
                
                r_data[15630] <= r_data[15629];
                
                r_data[15631] <= r_data[15630];
                
                r_data[15632] <= r_data[15631];
                
                r_data[15633] <= r_data[15632];
                
                r_data[15634] <= r_data[15633];
                
                r_data[15635] <= r_data[15634];
                
                r_data[15636] <= r_data[15635];
                
                r_data[15637] <= r_data[15636];
                
                r_data[15638] <= r_data[15637];
                
                r_data[15639] <= r_data[15638];
                
                r_data[15640] <= r_data[15639];
                
                r_data[15641] <= r_data[15640];
                
                r_data[15642] <= r_data[15641];
                
                r_data[15643] <= r_data[15642];
                
                r_data[15644] <= r_data[15643];
                
                r_data[15645] <= r_data[15644];
                
                r_data[15646] <= r_data[15645];
                
                r_data[15647] <= r_data[15646];
                
                r_data[15648] <= r_data[15647];
                
                r_data[15649] <= r_data[15648];
                
                r_data[15650] <= r_data[15649];
                
                r_data[15651] <= r_data[15650];
                
                r_data[15652] <= r_data[15651];
                
                r_data[15653] <= r_data[15652];
                
                r_data[15654] <= r_data[15653];
                
                r_data[15655] <= r_data[15654];
                
                r_data[15656] <= r_data[15655];
                
                r_data[15657] <= r_data[15656];
                
                r_data[15658] <= r_data[15657];
                
                r_data[15659] <= r_data[15658];
                
                r_data[15660] <= r_data[15659];
                
                r_data[15661] <= r_data[15660];
                
                r_data[15662] <= r_data[15661];
                
                r_data[15663] <= r_data[15662];
                
                r_data[15664] <= r_data[15663];
                
                r_data[15665] <= r_data[15664];
                
                r_data[15666] <= r_data[15665];
                
                r_data[15667] <= r_data[15666];
                
                r_data[15668] <= r_data[15667];
                
                r_data[15669] <= r_data[15668];
                
                r_data[15670] <= r_data[15669];
                
                r_data[15671] <= r_data[15670];
                
                r_data[15672] <= r_data[15671];
                
                r_data[15673] <= r_data[15672];
                
                r_data[15674] <= r_data[15673];
                
                r_data[15675] <= r_data[15674];
                
                r_data[15676] <= r_data[15675];
                
                r_data[15677] <= r_data[15676];
                
                r_data[15678] <= r_data[15677];
                
                r_data[15679] <= r_data[15678];
                
                r_data[15680] <= r_data[15679];
                
                r_data[15681] <= r_data[15680];
                
                r_data[15682] <= r_data[15681];
                
                r_data[15683] <= r_data[15682];
                
                r_data[15684] <= r_data[15683];
                
                r_data[15685] <= r_data[15684];
                
                r_data[15686] <= r_data[15685];
                
                r_data[15687] <= r_data[15686];
                
                r_data[15688] <= r_data[15687];
                
                r_data[15689] <= r_data[15688];
                
                r_data[15690] <= r_data[15689];
                
                r_data[15691] <= r_data[15690];
                
                r_data[15692] <= r_data[15691];
                
                r_data[15693] <= r_data[15692];
                
                r_data[15694] <= r_data[15693];
                
                r_data[15695] <= r_data[15694];
                
                r_data[15696] <= r_data[15695];
                
                r_data[15697] <= r_data[15696];
                
                r_data[15698] <= r_data[15697];
                
                r_data[15699] <= r_data[15698];
                
                r_data[15700] <= r_data[15699];
                
                r_data[15701] <= r_data[15700];
                
                r_data[15702] <= r_data[15701];
                
                r_data[15703] <= r_data[15702];
                
                r_data[15704] <= r_data[15703];
                
                r_data[15705] <= r_data[15704];
                
                r_data[15706] <= r_data[15705];
                
                r_data[15707] <= r_data[15706];
                
                r_data[15708] <= r_data[15707];
                
                r_data[15709] <= r_data[15708];
                
                r_data[15710] <= r_data[15709];
                
                r_data[15711] <= r_data[15710];
                
                r_data[15712] <= r_data[15711];
                
                r_data[15713] <= r_data[15712];
                
                r_data[15714] <= r_data[15713];
                
                r_data[15715] <= r_data[15714];
                
                r_data[15716] <= r_data[15715];
                
                r_data[15717] <= r_data[15716];
                
                r_data[15718] <= r_data[15717];
                
                r_data[15719] <= r_data[15718];
                
                r_data[15720] <= r_data[15719];
                
                r_data[15721] <= r_data[15720];
                
                r_data[15722] <= r_data[15721];
                
                r_data[15723] <= r_data[15722];
                
                r_data[15724] <= r_data[15723];
                
                r_data[15725] <= r_data[15724];
                
                r_data[15726] <= r_data[15725];
                
                r_data[15727] <= r_data[15726];
                
                r_data[15728] <= r_data[15727];
                
                r_data[15729] <= r_data[15728];
                
                r_data[15730] <= r_data[15729];
                
                r_data[15731] <= r_data[15730];
                
                r_data[15732] <= r_data[15731];
                
                r_data[15733] <= r_data[15732];
                
                r_data[15734] <= r_data[15733];
                
                r_data[15735] <= r_data[15734];
                
                r_data[15736] <= r_data[15735];
                
                r_data[15737] <= r_data[15736];
                
                r_data[15738] <= r_data[15737];
                
                r_data[15739] <= r_data[15738];
                
                r_data[15740] <= r_data[15739];
                
                r_data[15741] <= r_data[15740];
                
                r_data[15742] <= r_data[15741];
                
                r_data[15743] <= r_data[15742];
                
                r_data[15744] <= r_data[15743];
                
                r_data[15745] <= r_data[15744];
                
                r_data[15746] <= r_data[15745];
                
                r_data[15747] <= r_data[15746];
                
                r_data[15748] <= r_data[15747];
                
                r_data[15749] <= r_data[15748];
                
                r_data[15750] <= r_data[15749];
                
                r_data[15751] <= r_data[15750];
                
                r_data[15752] <= r_data[15751];
                
                r_data[15753] <= r_data[15752];
                
                r_data[15754] <= r_data[15753];
                
                r_data[15755] <= r_data[15754];
                
                r_data[15756] <= r_data[15755];
                
                r_data[15757] <= r_data[15756];
                
                r_data[15758] <= r_data[15757];
                
                r_data[15759] <= r_data[15758];
                
                r_data[15760] <= r_data[15759];
                
                r_data[15761] <= r_data[15760];
                
                r_data[15762] <= r_data[15761];
                
                r_data[15763] <= r_data[15762];
                
                r_data[15764] <= r_data[15763];
                
                r_data[15765] <= r_data[15764];
                
                r_data[15766] <= r_data[15765];
                
                r_data[15767] <= r_data[15766];
                
                r_data[15768] <= r_data[15767];
                
                r_data[15769] <= r_data[15768];
                
                r_data[15770] <= r_data[15769];
                
                r_data[15771] <= r_data[15770];
                
                r_data[15772] <= r_data[15771];
                
                r_data[15773] <= r_data[15772];
                
                r_data[15774] <= r_data[15773];
                
                r_data[15775] <= r_data[15774];
                
                r_data[15776] <= r_data[15775];
                
                r_data[15777] <= r_data[15776];
                
                r_data[15778] <= r_data[15777];
                
                r_data[15779] <= r_data[15778];
                
                r_data[15780] <= r_data[15779];
                
                r_data[15781] <= r_data[15780];
                
                r_data[15782] <= r_data[15781];
                
                r_data[15783] <= r_data[15782];
                
                r_data[15784] <= r_data[15783];
                
                r_data[15785] <= r_data[15784];
                
                r_data[15786] <= r_data[15785];
                
                r_data[15787] <= r_data[15786];
                
                r_data[15788] <= r_data[15787];
                
                r_data[15789] <= r_data[15788];
                
                r_data[15790] <= r_data[15789];
                
                r_data[15791] <= r_data[15790];
                
                r_data[15792] <= r_data[15791];
                
                r_data[15793] <= r_data[15792];
                
                r_data[15794] <= r_data[15793];
                
                r_data[15795] <= r_data[15794];
                
                r_data[15796] <= r_data[15795];
                
                r_data[15797] <= r_data[15796];
                
                r_data[15798] <= r_data[15797];
                
                r_data[15799] <= r_data[15798];
                
                r_data[15800] <= r_data[15799];
                
                r_data[15801] <= r_data[15800];
                
                r_data[15802] <= r_data[15801];
                
                r_data[15803] <= r_data[15802];
                
                r_data[15804] <= r_data[15803];
                
                r_data[15805] <= r_data[15804];
                
                r_data[15806] <= r_data[15805];
                
                r_data[15807] <= r_data[15806];
                
                r_data[15808] <= r_data[15807];
                
                r_data[15809] <= r_data[15808];
                
                r_data[15810] <= r_data[15809];
                
                r_data[15811] <= r_data[15810];
                
                r_data[15812] <= r_data[15811];
                
                r_data[15813] <= r_data[15812];
                
                r_data[15814] <= r_data[15813];
                
                r_data[15815] <= r_data[15814];
                
                r_data[15816] <= r_data[15815];
                
                r_data[15817] <= r_data[15816];
                
                r_data[15818] <= r_data[15817];
                
                r_data[15819] <= r_data[15818];
                
                r_data[15820] <= r_data[15819];
                
                r_data[15821] <= r_data[15820];
                
                r_data[15822] <= r_data[15821];
                
                r_data[15823] <= r_data[15822];
                
                r_data[15824] <= r_data[15823];
                
                r_data[15825] <= r_data[15824];
                
                r_data[15826] <= r_data[15825];
                
                r_data[15827] <= r_data[15826];
                
                r_data[15828] <= r_data[15827];
                
                r_data[15829] <= r_data[15828];
                
                r_data[15830] <= r_data[15829];
                
                r_data[15831] <= r_data[15830];
                
                r_data[15832] <= r_data[15831];
                
                r_data[15833] <= r_data[15832];
                
                r_data[15834] <= r_data[15833];
                
                r_data[15835] <= r_data[15834];
                
                r_data[15836] <= r_data[15835];
                
                r_data[15837] <= r_data[15836];
                
                r_data[15838] <= r_data[15837];
                
                r_data[15839] <= r_data[15838];
                
                r_data[15840] <= r_data[15839];
                
                r_data[15841] <= r_data[15840];
                
                r_data[15842] <= r_data[15841];
                
                r_data[15843] <= r_data[15842];
                
                r_data[15844] <= r_data[15843];
                
                r_data[15845] <= r_data[15844];
                
                r_data[15846] <= r_data[15845];
                
                r_data[15847] <= r_data[15846];
                
                r_data[15848] <= r_data[15847];
                
                r_data[15849] <= r_data[15848];
                
                r_data[15850] <= r_data[15849];
                
                r_data[15851] <= r_data[15850];
                
                r_data[15852] <= r_data[15851];
                
                r_data[15853] <= r_data[15852];
                
                r_data[15854] <= r_data[15853];
                
                r_data[15855] <= r_data[15854];
                
                r_data[15856] <= r_data[15855];
                
                r_data[15857] <= r_data[15856];
                
                r_data[15858] <= r_data[15857];
                
                r_data[15859] <= r_data[15858];
                
                r_data[15860] <= r_data[15859];
                
                r_data[15861] <= r_data[15860];
                
                r_data[15862] <= r_data[15861];
                
                r_data[15863] <= r_data[15862];
                
                r_data[15864] <= r_data[15863];
                
                r_data[15865] <= r_data[15864];
                
                r_data[15866] <= r_data[15865];
                
                r_data[15867] <= r_data[15866];
                
                r_data[15868] <= r_data[15867];
                
                r_data[15869] <= r_data[15868];
                
                r_data[15870] <= r_data[15869];
                
                r_data[15871] <= r_data[15870];
                
                r_data[15872] <= r_data[15871];
                
                r_data[15873] <= r_data[15872];
                
                r_data[15874] <= r_data[15873];
                
                r_data[15875] <= r_data[15874];
                
                r_data[15876] <= r_data[15875];
                
                r_data[15877] <= r_data[15876];
                
                r_data[15878] <= r_data[15877];
                
                r_data[15879] <= r_data[15878];
                
                r_data[15880] <= r_data[15879];
                
                r_data[15881] <= r_data[15880];
                
                r_data[15882] <= r_data[15881];
                
                r_data[15883] <= r_data[15882];
                
                r_data[15884] <= r_data[15883];
                
                r_data[15885] <= r_data[15884];
                
                r_data[15886] <= r_data[15885];
                
                r_data[15887] <= r_data[15886];
                
                r_data[15888] <= r_data[15887];
                
                r_data[15889] <= r_data[15888];
                
                r_data[15890] <= r_data[15889];
                
                r_data[15891] <= r_data[15890];
                
                r_data[15892] <= r_data[15891];
                
                r_data[15893] <= r_data[15892];
                
                r_data[15894] <= r_data[15893];
                
                r_data[15895] <= r_data[15894];
                
                r_data[15896] <= r_data[15895];
                
                r_data[15897] <= r_data[15896];
                
                r_data[15898] <= r_data[15897];
                
                r_data[15899] <= r_data[15898];
                
                r_data[15900] <= r_data[15899];
                
                r_data[15901] <= r_data[15900];
                
                r_data[15902] <= r_data[15901];
                
                r_data[15903] <= r_data[15902];
                
                r_data[15904] <= r_data[15903];
                
                r_data[15905] <= r_data[15904];
                
                r_data[15906] <= r_data[15905];
                
                r_data[15907] <= r_data[15906];
                
                r_data[15908] <= r_data[15907];
                
                r_data[15909] <= r_data[15908];
                
                r_data[15910] <= r_data[15909];
                
                r_data[15911] <= r_data[15910];
                
                r_data[15912] <= r_data[15911];
                
                r_data[15913] <= r_data[15912];
                
                r_data[15914] <= r_data[15913];
                
                r_data[15915] <= r_data[15914];
                
                r_data[15916] <= r_data[15915];
                
                r_data[15917] <= r_data[15916];
                
                r_data[15918] <= r_data[15917];
                
                r_data[15919] <= r_data[15918];
                
                r_data[15920] <= r_data[15919];
                
                r_data[15921] <= r_data[15920];
                
                r_data[15922] <= r_data[15921];
                
                r_data[15923] <= r_data[15922];
                
                r_data[15924] <= r_data[15923];
                
                r_data[15925] <= r_data[15924];
                
                r_data[15926] <= r_data[15925];
                
                r_data[15927] <= r_data[15926];
                
                r_data[15928] <= r_data[15927];
                
                r_data[15929] <= r_data[15928];
                
                r_data[15930] <= r_data[15929];
                
                r_data[15931] <= r_data[15930];
                
                r_data[15932] <= r_data[15931];
                
                r_data[15933] <= r_data[15932];
                
                r_data[15934] <= r_data[15933];
                
                r_data[15935] <= r_data[15934];
                
                r_data[15936] <= r_data[15935];
                
                r_data[15937] <= r_data[15936];
                
                r_data[15938] <= r_data[15937];
                
                r_data[15939] <= r_data[15938];
                
                r_data[15940] <= r_data[15939];
                
                r_data[15941] <= r_data[15940];
                
                r_data[15942] <= r_data[15941];
                
                r_data[15943] <= r_data[15942];
                
                r_data[15944] <= r_data[15943];
                
                r_data[15945] <= r_data[15944];
                
                r_data[15946] <= r_data[15945];
                
                r_data[15947] <= r_data[15946];
                
                r_data[15948] <= r_data[15947];
                
                r_data[15949] <= r_data[15948];
                
                r_data[15950] <= r_data[15949];
                
                r_data[15951] <= r_data[15950];
                
                r_data[15952] <= r_data[15951];
                
                r_data[15953] <= r_data[15952];
                
                r_data[15954] <= r_data[15953];
                
                r_data[15955] <= r_data[15954];
                
                r_data[15956] <= r_data[15955];
                
                r_data[15957] <= r_data[15956];
                
                r_data[15958] <= r_data[15957];
                
                r_data[15959] <= r_data[15958];
                
                r_data[15960] <= r_data[15959];
                
                r_data[15961] <= r_data[15960];
                
                r_data[15962] <= r_data[15961];
                
                r_data[15963] <= r_data[15962];
                
                r_data[15964] <= r_data[15963];
                
                r_data[15965] <= r_data[15964];
                
                r_data[15966] <= r_data[15965];
                
                r_data[15967] <= r_data[15966];
                
                r_data[15968] <= r_data[15967];
                
                r_data[15969] <= r_data[15968];
                
                r_data[15970] <= r_data[15969];
                
                r_data[15971] <= r_data[15970];
                
                r_data[15972] <= r_data[15971];
                
                r_data[15973] <= r_data[15972];
                
                r_data[15974] <= r_data[15973];
                
                r_data[15975] <= r_data[15974];
                
                r_data[15976] <= r_data[15975];
                
                r_data[15977] <= r_data[15976];
                
                r_data[15978] <= r_data[15977];
                
                r_data[15979] <= r_data[15978];
                
                r_data[15980] <= r_data[15979];
                
                r_data[15981] <= r_data[15980];
                
                r_data[15982] <= r_data[15981];
                
                r_data[15983] <= r_data[15982];
                
                r_data[15984] <= r_data[15983];
                
                r_data[15985] <= r_data[15984];
                
                r_data[15986] <= r_data[15985];
                
                r_data[15987] <= r_data[15986];
                
                r_data[15988] <= r_data[15987];
                
                r_data[15989] <= r_data[15988];
                
                r_data[15990] <= r_data[15989];
                
                r_data[15991] <= r_data[15990];
                
                r_data[15992] <= r_data[15991];
                
                r_data[15993] <= r_data[15992];
                
                r_data[15994] <= r_data[15993];
                
                r_data[15995] <= r_data[15994];
                
                r_data[15996] <= r_data[15995];
                
                r_data[15997] <= r_data[15996];
                
                r_data[15998] <= r_data[15997];
                
                r_data[15999] <= r_data[15998];
                
                r_data[16000] <= r_data[15999];
                
                r_data[16001] <= r_data[16000];
                
                r_data[16002] <= r_data[16001];
                
                r_data[16003] <= r_data[16002];
                
                r_data[16004] <= r_data[16003];
                
                r_data[16005] <= r_data[16004];
                
                r_data[16006] <= r_data[16005];
                
                r_data[16007] <= r_data[16006];
                
                r_data[16008] <= r_data[16007];
                
                r_data[16009] <= r_data[16008];
                
                r_data[16010] <= r_data[16009];
                
                r_data[16011] <= r_data[16010];
                
                r_data[16012] <= r_data[16011];
                
                r_data[16013] <= r_data[16012];
                
                r_data[16014] <= r_data[16013];
                
                r_data[16015] <= r_data[16014];
                
                r_data[16016] <= r_data[16015];
                
                r_data[16017] <= r_data[16016];
                
                r_data[16018] <= r_data[16017];
                
                r_data[16019] <= r_data[16018];
                
                r_data[16020] <= r_data[16019];
                
                r_data[16021] <= r_data[16020];
                
                r_data[16022] <= r_data[16021];
                
                r_data[16023] <= r_data[16022];
                
                r_data[16024] <= r_data[16023];
                
                r_data[16025] <= r_data[16024];
                
                r_data[16026] <= r_data[16025];
                
                r_data[16027] <= r_data[16026];
                
                r_data[16028] <= r_data[16027];
                
                r_data[16029] <= r_data[16028];
                
                r_data[16030] <= r_data[16029];
                
                r_data[16031] <= r_data[16030];
                
                r_data[16032] <= r_data[16031];
                
                r_data[16033] <= r_data[16032];
                
                r_data[16034] <= r_data[16033];
                
                r_data[16035] <= r_data[16034];
                
                r_data[16036] <= r_data[16035];
                
                r_data[16037] <= r_data[16036];
                
                r_data[16038] <= r_data[16037];
                
                r_data[16039] <= r_data[16038];
                
                r_data[16040] <= r_data[16039];
                
                r_data[16041] <= r_data[16040];
                
                r_data[16042] <= r_data[16041];
                
                r_data[16043] <= r_data[16042];
                
                r_data[16044] <= r_data[16043];
                
                r_data[16045] <= r_data[16044];
                
                r_data[16046] <= r_data[16045];
                
                r_data[16047] <= r_data[16046];
                
                r_data[16048] <= r_data[16047];
                
                r_data[16049] <= r_data[16048];
                
                r_data[16050] <= r_data[16049];
                
                r_data[16051] <= r_data[16050];
                
                r_data[16052] <= r_data[16051];
                
                r_data[16053] <= r_data[16052];
                
                r_data[16054] <= r_data[16053];
                
                r_data[16055] <= r_data[16054];
                
                r_data[16056] <= r_data[16055];
                
                r_data[16057] <= r_data[16056];
                
                r_data[16058] <= r_data[16057];
                
                r_data[16059] <= r_data[16058];
                
                r_data[16060] <= r_data[16059];
                
                r_data[16061] <= r_data[16060];
                
                r_data[16062] <= r_data[16061];
                
                r_data[16063] <= r_data[16062];
                
                r_data[16064] <= r_data[16063];
                
                r_data[16065] <= r_data[16064];
                
                r_data[16066] <= r_data[16065];
                
                r_data[16067] <= r_data[16066];
                
                r_data[16068] <= r_data[16067];
                
                r_data[16069] <= r_data[16068];
                
                r_data[16070] <= r_data[16069];
                
                r_data[16071] <= r_data[16070];
                
                r_data[16072] <= r_data[16071];
                
                r_data[16073] <= r_data[16072];
                
                r_data[16074] <= r_data[16073];
                
                r_data[16075] <= r_data[16074];
                
                r_data[16076] <= r_data[16075];
                
                r_data[16077] <= r_data[16076];
                
                r_data[16078] <= r_data[16077];
                
                r_data[16079] <= r_data[16078];
                
                r_data[16080] <= r_data[16079];
                
                r_data[16081] <= r_data[16080];
                
                r_data[16082] <= r_data[16081];
                
                r_data[16083] <= r_data[16082];
                
                r_data[16084] <= r_data[16083];
                
                r_data[16085] <= r_data[16084];
                
                r_data[16086] <= r_data[16085];
                
                r_data[16087] <= r_data[16086];
                
                r_data[16088] <= r_data[16087];
                
                r_data[16089] <= r_data[16088];
                
                r_data[16090] <= r_data[16089];
                
                r_data[16091] <= r_data[16090];
                
                r_data[16092] <= r_data[16091];
                
                r_data[16093] <= r_data[16092];
                
                r_data[16094] <= r_data[16093];
                
                r_data[16095] <= r_data[16094];
                
                r_data[16096] <= r_data[16095];
                
                r_data[16097] <= r_data[16096];
                
                r_data[16098] <= r_data[16097];
                
                r_data[16099] <= r_data[16098];
                
                r_data[16100] <= r_data[16099];
                
                r_data[16101] <= r_data[16100];
                
                r_data[16102] <= r_data[16101];
                
                r_data[16103] <= r_data[16102];
                
                r_data[16104] <= r_data[16103];
                
                r_data[16105] <= r_data[16104];
                
                r_data[16106] <= r_data[16105];
                
                r_data[16107] <= r_data[16106];
                
                r_data[16108] <= r_data[16107];
                
                r_data[16109] <= r_data[16108];
                
                r_data[16110] <= r_data[16109];
                
                r_data[16111] <= r_data[16110];
                
                r_data[16112] <= r_data[16111];
                
                r_data[16113] <= r_data[16112];
                
                r_data[16114] <= r_data[16113];
                
                r_data[16115] <= r_data[16114];
                
                r_data[16116] <= r_data[16115];
                
                r_data[16117] <= r_data[16116];
                
                r_data[16118] <= r_data[16117];
                
                r_data[16119] <= r_data[16118];
                
                r_data[16120] <= r_data[16119];
                
                r_data[16121] <= r_data[16120];
                
                r_data[16122] <= r_data[16121];
                
                r_data[16123] <= r_data[16122];
                
                r_data[16124] <= r_data[16123];
                
                r_data[16125] <= r_data[16124];
                
                r_data[16126] <= r_data[16125];
                
                r_data[16127] <= r_data[16126];
                
                r_data[16128] <= r_data[16127];
                
                r_data[16129] <= r_data[16128];
                
                r_data[16130] <= r_data[16129];
                
                r_data[16131] <= r_data[16130];
                
                r_data[16132] <= r_data[16131];
                
                r_data[16133] <= r_data[16132];
                
                r_data[16134] <= r_data[16133];
                
                r_data[16135] <= r_data[16134];
                
                r_data[16136] <= r_data[16135];
                
                r_data[16137] <= r_data[16136];
                
                r_data[16138] <= r_data[16137];
                
                r_data[16139] <= r_data[16138];
                
                r_data[16140] <= r_data[16139];
                
                r_data[16141] <= r_data[16140];
                
                r_data[16142] <= r_data[16141];
                
                r_data[16143] <= r_data[16142];
                
                r_data[16144] <= r_data[16143];
                
                r_data[16145] <= r_data[16144];
                
                r_data[16146] <= r_data[16145];
                
                r_data[16147] <= r_data[16146];
                
                r_data[16148] <= r_data[16147];
                
                r_data[16149] <= r_data[16148];
                
                r_data[16150] <= r_data[16149];
                
                r_data[16151] <= r_data[16150];
                
                r_data[16152] <= r_data[16151];
                
                r_data[16153] <= r_data[16152];
                
                r_data[16154] <= r_data[16153];
                
                r_data[16155] <= r_data[16154];
                
                r_data[16156] <= r_data[16155];
                
                r_data[16157] <= r_data[16156];
                
                r_data[16158] <= r_data[16157];
                
                r_data[16159] <= r_data[16158];
                
                r_data[16160] <= r_data[16159];
                
                r_data[16161] <= r_data[16160];
                
                r_data[16162] <= r_data[16161];
                
                r_data[16163] <= r_data[16162];
                
                r_data[16164] <= r_data[16163];
                
                r_data[16165] <= r_data[16164];
                
                r_data[16166] <= r_data[16165];
                
                r_data[16167] <= r_data[16166];
                
                r_data[16168] <= r_data[16167];
                
                r_data[16169] <= r_data[16168];
                
                r_data[16170] <= r_data[16169];
                
                r_data[16171] <= r_data[16170];
                
                r_data[16172] <= r_data[16171];
                
                r_data[16173] <= r_data[16172];
                
                r_data[16174] <= r_data[16173];
                
                r_data[16175] <= r_data[16174];
                
                r_data[16176] <= r_data[16175];
                
                r_data[16177] <= r_data[16176];
                
                r_data[16178] <= r_data[16177];
                
                r_data[16179] <= r_data[16178];
                
                r_data[16180] <= r_data[16179];
                
                r_data[16181] <= r_data[16180];
                
                r_data[16182] <= r_data[16181];
                
                r_data[16183] <= r_data[16182];
                
                r_data[16184] <= r_data[16183];
                
                r_data[16185] <= r_data[16184];
                
                r_data[16186] <= r_data[16185];
                
                r_data[16187] <= r_data[16186];
                
                r_data[16188] <= r_data[16187];
                
                r_data[16189] <= r_data[16188];
                
                r_data[16190] <= r_data[16189];
                
                r_data[16191] <= r_data[16190];
                
                r_data[16192] <= r_data[16191];
                
                r_data[16193] <= r_data[16192];
                
                r_data[16194] <= r_data[16193];
                
                r_data[16195] <= r_data[16194];
                
                r_data[16196] <= r_data[16195];
                
                r_data[16197] <= r_data[16196];
                
                r_data[16198] <= r_data[16197];
                
                r_data[16199] <= r_data[16198];
                
                r_data[16200] <= r_data[16199];
                
                r_data[16201] <= r_data[16200];
                
                r_data[16202] <= r_data[16201];
                
                r_data[16203] <= r_data[16202];
                
                r_data[16204] <= r_data[16203];
                
                r_data[16205] <= r_data[16204];
                
                r_data[16206] <= r_data[16205];
                
                r_data[16207] <= r_data[16206];
                
                r_data[16208] <= r_data[16207];
                
                r_data[16209] <= r_data[16208];
                
                r_data[16210] <= r_data[16209];
                
                r_data[16211] <= r_data[16210];
                
                r_data[16212] <= r_data[16211];
                
                r_data[16213] <= r_data[16212];
                
                r_data[16214] <= r_data[16213];
                
                r_data[16215] <= r_data[16214];
                
                r_data[16216] <= r_data[16215];
                
                r_data[16217] <= r_data[16216];
                
                r_data[16218] <= r_data[16217];
                
                r_data[16219] <= r_data[16218];
                
                r_data[16220] <= r_data[16219];
                
                r_data[16221] <= r_data[16220];
                
                r_data[16222] <= r_data[16221];
                
                r_data[16223] <= r_data[16222];
                
                r_data[16224] <= r_data[16223];
                
                r_data[16225] <= r_data[16224];
                
                r_data[16226] <= r_data[16225];
                
                r_data[16227] <= r_data[16226];
                
                r_data[16228] <= r_data[16227];
                
                r_data[16229] <= r_data[16228];
                
                r_data[16230] <= r_data[16229];
                
                r_data[16231] <= r_data[16230];
                
                r_data[16232] <= r_data[16231];
                
                r_data[16233] <= r_data[16232];
                
                r_data[16234] <= r_data[16233];
                
                r_data[16235] <= r_data[16234];
                
                r_data[16236] <= r_data[16235];
                
                r_data[16237] <= r_data[16236];
                
                r_data[16238] <= r_data[16237];
                
                r_data[16239] <= r_data[16238];
                
                r_data[16240] <= r_data[16239];
                
                r_data[16241] <= r_data[16240];
                
                r_data[16242] <= r_data[16241];
                
                r_data[16243] <= r_data[16242];
                
                r_data[16244] <= r_data[16243];
                
                r_data[16245] <= r_data[16244];
                
                r_data[16246] <= r_data[16245];
                
                r_data[16247] <= r_data[16246];
                
                r_data[16248] <= r_data[16247];
                
                r_data[16249] <= r_data[16248];
                
                r_data[16250] <= r_data[16249];
                
                r_data[16251] <= r_data[16250];
                
                r_data[16252] <= r_data[16251];
                
                r_data[16253] <= r_data[16252];
                
                r_data[16254] <= r_data[16253];
                
                r_data[16255] <= r_data[16254];
                
                r_data[16256] <= r_data[16255];
                
                r_data[16257] <= r_data[16256];
                
                r_data[16258] <= r_data[16257];
                
                r_data[16259] <= r_data[16258];
                
                r_data[16260] <= r_data[16259];
                
                r_data[16261] <= r_data[16260];
                
                r_data[16262] <= r_data[16261];
                
                r_data[16263] <= r_data[16262];
                
                r_data[16264] <= r_data[16263];
                
                r_data[16265] <= r_data[16264];
                
                r_data[16266] <= r_data[16265];
                
                r_data[16267] <= r_data[16266];
                
                r_data[16268] <= r_data[16267];
                
                r_data[16269] <= r_data[16268];
                
                r_data[16270] <= r_data[16269];
                
                r_data[16271] <= r_data[16270];
                
                r_data[16272] <= r_data[16271];
                
                r_data[16273] <= r_data[16272];
                
                r_data[16274] <= r_data[16273];
                
                r_data[16275] <= r_data[16274];
                
                r_data[16276] <= r_data[16275];
                
                r_data[16277] <= r_data[16276];
                
                r_data[16278] <= r_data[16277];
                
                r_data[16279] <= r_data[16278];
                
                r_data[16280] <= r_data[16279];
                
                r_data[16281] <= r_data[16280];
                
                r_data[16282] <= r_data[16281];
                
                r_data[16283] <= r_data[16282];
                
                r_data[16284] <= r_data[16283];
                
                r_data[16285] <= r_data[16284];
                
                r_data[16286] <= r_data[16285];
                
                r_data[16287] <= r_data[16286];
                
                r_data[16288] <= r_data[16287];
                
                r_data[16289] <= r_data[16288];
                
                r_data[16290] <= r_data[16289];
                
                r_data[16291] <= r_data[16290];
                
                r_data[16292] <= r_data[16291];
                
                r_data[16293] <= r_data[16292];
                
                r_data[16294] <= r_data[16293];
                
                r_data[16295] <= r_data[16294];
                
                r_data[16296] <= r_data[16295];
                
                r_data[16297] <= r_data[16296];
                
                r_data[16298] <= r_data[16297];
                
                r_data[16299] <= r_data[16298];
                
                r_data[16300] <= r_data[16299];
                
                r_data[16301] <= r_data[16300];
                
                r_data[16302] <= r_data[16301];
                
                r_data[16303] <= r_data[16302];
                
                r_data[16304] <= r_data[16303];
                
                r_data[16305] <= r_data[16304];
                
                r_data[16306] <= r_data[16305];
                
                r_data[16307] <= r_data[16306];
                
                r_data[16308] <= r_data[16307];
                
                r_data[16309] <= r_data[16308];
                
                r_data[16310] <= r_data[16309];
                
                r_data[16311] <= r_data[16310];
                
                r_data[16312] <= r_data[16311];
                
                r_data[16313] <= r_data[16312];
                
                r_data[16314] <= r_data[16313];
                
                r_data[16315] <= r_data[16314];
                
                r_data[16316] <= r_data[16315];
                
                r_data[16317] <= r_data[16316];
                
                r_data[16318] <= r_data[16317];
                
                r_data[16319] <= r_data[16318];
                
                r_data[16320] <= r_data[16319];
                
                r_data[16321] <= r_data[16320];
                
                r_data[16322] <= r_data[16321];
                
                r_data[16323] <= r_data[16322];
                
                r_data[16324] <= r_data[16323];
                
                r_data[16325] <= r_data[16324];
                
                r_data[16326] <= r_data[16325];
                
                r_data[16327] <= r_data[16326];
                
                r_data[16328] <= r_data[16327];
                
                r_data[16329] <= r_data[16328];
                
                r_data[16330] <= r_data[16329];
                
                r_data[16331] <= r_data[16330];
                
                r_data[16332] <= r_data[16331];
                
                r_data[16333] <= r_data[16332];
                
                r_data[16334] <= r_data[16333];
                
                r_data[16335] <= r_data[16334];
                
                r_data[16336] <= r_data[16335];
                
                r_data[16337] <= r_data[16336];
                
                r_data[16338] <= r_data[16337];
                
                r_data[16339] <= r_data[16338];
                
                r_data[16340] <= r_data[16339];
                
                r_data[16341] <= r_data[16340];
                
                r_data[16342] <= r_data[16341];
                
                r_data[16343] <= r_data[16342];
                
                r_data[16344] <= r_data[16343];
                
                r_data[16345] <= r_data[16344];
                
                r_data[16346] <= r_data[16345];
                
                r_data[16347] <= r_data[16346];
                
                r_data[16348] <= r_data[16347];
                
                r_data[16349] <= r_data[16348];
                
                r_data[16350] <= r_data[16349];
                
                r_data[16351] <= r_data[16350];
                
                r_data[16352] <= r_data[16351];
                
                r_data[16353] <= r_data[16352];
                
                r_data[16354] <= r_data[16353];
                
                r_data[16355] <= r_data[16354];
                
                r_data[16356] <= r_data[16355];
                
                r_data[16357] <= r_data[16356];
                
                r_data[16358] <= r_data[16357];
                
                r_data[16359] <= r_data[16358];
                
                r_data[16360] <= r_data[16359];
                
                r_data[16361] <= r_data[16360];
                
                r_data[16362] <= r_data[16361];
                
                r_data[16363] <= r_data[16362];
                
                r_data[16364] <= r_data[16363];
                
                r_data[16365] <= r_data[16364];
                
                r_data[16366] <= r_data[16365];
                
                r_data[16367] <= r_data[16366];
                
                r_data[16368] <= r_data[16367];
                
                r_data[16369] <= r_data[16368];
                
                r_data[16370] <= r_data[16369];
                
                r_data[16371] <= r_data[16370];
                
                r_data[16372] <= r_data[16371];
                
                r_data[16373] <= r_data[16372];
                
                r_data[16374] <= r_data[16373];
                
                r_data[16375] <= r_data[16374];
                
                r_data[16376] <= r_data[16375];
                
                r_data[16377] <= r_data[16376];
                
                r_data[16378] <= r_data[16377];
                
                r_data[16379] <= r_data[16378];
                
                r_data[16380] <= r_data[16379];
                
                r_data[16381] <= r_data[16380];
                
                r_data[16382] <= r_data[16381];
                
                r_data[16383] <= r_data[16382];
                
                r_data[16384] <= r_data[16383];
                
                r_data[16385] <= r_data[16384];
                
                r_data[16386] <= r_data[16385];
                
                r_data[16387] <= r_data[16386];
                
                r_data[16388] <= r_data[16387];
                
                r_data[16389] <= r_data[16388];
                
                r_data[16390] <= r_data[16389];
                
                r_data[16391] <= r_data[16390];
                
                r_data[16392] <= r_data[16391];
                
                r_data[16393] <= r_data[16392];
                
                r_data[16394] <= r_data[16393];
                
                r_data[16395] <= r_data[16394];
                
                r_data[16396] <= r_data[16395];
                
                r_data[16397] <= r_data[16396];
                
                r_data[16398] <= r_data[16397];
                
                r_data[16399] <= r_data[16398];
                
                r_data[16400] <= r_data[16399];
                
                r_data[16401] <= r_data[16400];
                
                r_data[16402] <= r_data[16401];
                
                r_data[16403] <= r_data[16402];
                
                r_data[16404] <= r_data[16403];
                
                r_data[16405] <= r_data[16404];
                
                r_data[16406] <= r_data[16405];
                
                r_data[16407] <= r_data[16406];
                
                r_data[16408] <= r_data[16407];
                
                r_data[16409] <= r_data[16408];
                
                r_data[16410] <= r_data[16409];
                
                r_data[16411] <= r_data[16410];
                
                r_data[16412] <= r_data[16411];
                
                r_data[16413] <= r_data[16412];
                
                r_data[16414] <= r_data[16413];
                
                r_data[16415] <= r_data[16414];
                
                r_data[16416] <= r_data[16415];
                
                r_data[16417] <= r_data[16416];
                
                r_data[16418] <= r_data[16417];
                
                r_data[16419] <= r_data[16418];
                
                r_data[16420] <= r_data[16419];
                
                r_data[16421] <= r_data[16420];
                
                r_data[16422] <= r_data[16421];
                
                r_data[16423] <= r_data[16422];
                
                r_data[16424] <= r_data[16423];
                
                r_data[16425] <= r_data[16424];
                
                r_data[16426] <= r_data[16425];
                
                r_data[16427] <= r_data[16426];
                
                r_data[16428] <= r_data[16427];
                
                r_data[16429] <= r_data[16428];
                
                r_data[16430] <= r_data[16429];
                
                r_data[16431] <= r_data[16430];
                
                r_data[16432] <= r_data[16431];
                
                r_data[16433] <= r_data[16432];
                
                r_data[16434] <= r_data[16433];
                
                r_data[16435] <= r_data[16434];
                
                r_data[16436] <= r_data[16435];
                
                r_data[16437] <= r_data[16436];
                
                r_data[16438] <= r_data[16437];
                
                r_data[16439] <= r_data[16438];
                
                r_data[16440] <= r_data[16439];
                
                r_data[16441] <= r_data[16440];
                
                r_data[16442] <= r_data[16441];
                
                r_data[16443] <= r_data[16442];
                
                r_data[16444] <= r_data[16443];
                
                r_data[16445] <= r_data[16444];
                
                r_data[16446] <= r_data[16445];
                
                r_data[16447] <= r_data[16446];
                
                r_data[16448] <= r_data[16447];
                
                r_data[16449] <= r_data[16448];
                
                r_data[16450] <= r_data[16449];
                
                r_data[16451] <= r_data[16450];
                
                r_data[16452] <= r_data[16451];
                
                r_data[16453] <= r_data[16452];
                
                r_data[16454] <= r_data[16453];
                
                r_data[16455] <= r_data[16454];
                
                r_data[16456] <= r_data[16455];
                
                r_data[16457] <= r_data[16456];
                
                r_data[16458] <= r_data[16457];
                
                r_data[16459] <= r_data[16458];
                
                r_data[16460] <= r_data[16459];
                
                r_data[16461] <= r_data[16460];
                
                r_data[16462] <= r_data[16461];
                
                r_data[16463] <= r_data[16462];
                
                r_data[16464] <= r_data[16463];
                
                r_data[16465] <= r_data[16464];
                
                r_data[16466] <= r_data[16465];
                
                r_data[16467] <= r_data[16466];
                
                r_data[16468] <= r_data[16467];
                
                r_data[16469] <= r_data[16468];
                
                r_data[16470] <= r_data[16469];
                
                r_data[16471] <= r_data[16470];
                
                r_data[16472] <= r_data[16471];
                
                r_data[16473] <= r_data[16472];
                
                r_data[16474] <= r_data[16473];
                
                r_data[16475] <= r_data[16474];
                
                r_data[16476] <= r_data[16475];
                
                r_data[16477] <= r_data[16476];
                
                r_data[16478] <= r_data[16477];
                
                r_data[16479] <= r_data[16478];
                
                r_data[16480] <= r_data[16479];
                
                r_data[16481] <= r_data[16480];
                
                r_data[16482] <= r_data[16481];
                
                r_data[16483] <= r_data[16482];
                
                r_data[16484] <= r_data[16483];
                
                r_data[16485] <= r_data[16484];
                
                r_data[16486] <= r_data[16485];
                
                r_data[16487] <= r_data[16486];
                
                r_data[16488] <= r_data[16487];
                
                r_data[16489] <= r_data[16488];
                
                r_data[16490] <= r_data[16489];
                
                r_data[16491] <= r_data[16490];
                
                r_data[16492] <= r_data[16491];
                
                r_data[16493] <= r_data[16492];
                
                r_data[16494] <= r_data[16493];
                
                r_data[16495] <= r_data[16494];
                
                r_data[16496] <= r_data[16495];
                
                r_data[16497] <= r_data[16496];
                
                r_data[16498] <= r_data[16497];
                
                r_data[16499] <= r_data[16498];
                
                r_data[16500] <= r_data[16499];
                
                r_data[16501] <= r_data[16500];
                
                r_data[16502] <= r_data[16501];
                
                r_data[16503] <= r_data[16502];
                
                r_data[16504] <= r_data[16503];
                
                r_data[16505] <= r_data[16504];
                
                r_data[16506] <= r_data[16505];
                
                r_data[16507] <= r_data[16506];
                
                r_data[16508] <= r_data[16507];
                
                r_data[16509] <= r_data[16508];
                
                r_data[16510] <= r_data[16509];
                
                r_data[16511] <= r_data[16510];
                
                r_data[16512] <= r_data[16511];
                
                r_data[16513] <= r_data[16512];
                
                r_data[16514] <= r_data[16513];
                
                r_data[16515] <= r_data[16514];
                
                r_data[16516] <= r_data[16515];
                
                r_data[16517] <= r_data[16516];
                
                r_data[16518] <= r_data[16517];
                
                r_data[16519] <= r_data[16518];
                
                r_data[16520] <= r_data[16519];
                
                r_data[16521] <= r_data[16520];
                
                r_data[16522] <= r_data[16521];
                
                r_data[16523] <= r_data[16522];
                
                r_data[16524] <= r_data[16523];
                
                r_data[16525] <= r_data[16524];
                
                r_data[16526] <= r_data[16525];
                
                r_data[16527] <= r_data[16526];
                
                r_data[16528] <= r_data[16527];
                
                r_data[16529] <= r_data[16528];
                
                r_data[16530] <= r_data[16529];
                
                r_data[16531] <= r_data[16530];
                
                r_data[16532] <= r_data[16531];
                
                r_data[16533] <= r_data[16532];
                
                r_data[16534] <= r_data[16533];
                
                r_data[16535] <= r_data[16534];
                
                r_data[16536] <= r_data[16535];
                
                r_data[16537] <= r_data[16536];
                
                r_data[16538] <= r_data[16537];
                
                r_data[16539] <= r_data[16538];
                
                r_data[16540] <= r_data[16539];
                
                r_data[16541] <= r_data[16540];
                
                r_data[16542] <= r_data[16541];
                
                r_data[16543] <= r_data[16542];
                
                r_data[16544] <= r_data[16543];
                
                r_data[16545] <= r_data[16544];
                
                r_data[16546] <= r_data[16545];
                
                r_data[16547] <= r_data[16546];
                
                r_data[16548] <= r_data[16547];
                
                r_data[16549] <= r_data[16548];
                
                r_data[16550] <= r_data[16549];
                
                r_data[16551] <= r_data[16550];
                
                r_data[16552] <= r_data[16551];
                
                r_data[16553] <= r_data[16552];
                
                r_data[16554] <= r_data[16553];
                
                r_data[16555] <= r_data[16554];
                
                r_data[16556] <= r_data[16555];
                
                r_data[16557] <= r_data[16556];
                
                r_data[16558] <= r_data[16557];
                
                r_data[16559] <= r_data[16558];
                
                r_data[16560] <= r_data[16559];
                
                r_data[16561] <= r_data[16560];
                
                r_data[16562] <= r_data[16561];
                
                r_data[16563] <= r_data[16562];
                
                r_data[16564] <= r_data[16563];
                
                r_data[16565] <= r_data[16564];
                
                r_data[16566] <= r_data[16565];
                
                r_data[16567] <= r_data[16566];
                
                r_data[16568] <= r_data[16567];
                
                r_data[16569] <= r_data[16568];
                
                r_data[16570] <= r_data[16569];
                
                r_data[16571] <= r_data[16570];
                
                r_data[16572] <= r_data[16571];
                
                r_data[16573] <= r_data[16572];
                
                r_data[16574] <= r_data[16573];
                
                r_data[16575] <= r_data[16574];
                
                r_data[16576] <= r_data[16575];
                
                r_data[16577] <= r_data[16576];
                
                r_data[16578] <= r_data[16577];
                
                r_data[16579] <= r_data[16578];
                
                r_data[16580] <= r_data[16579];
                
                r_data[16581] <= r_data[16580];
                
                r_data[16582] <= r_data[16581];
                
                r_data[16583] <= r_data[16582];
                
                r_data[16584] <= r_data[16583];
                
                r_data[16585] <= r_data[16584];
                
                r_data[16586] <= r_data[16585];
                
                r_data[16587] <= r_data[16586];
                
                r_data[16588] <= r_data[16587];
                
                r_data[16589] <= r_data[16588];
                
                r_data[16590] <= r_data[16589];
                
                r_data[16591] <= r_data[16590];
                
                r_data[16592] <= r_data[16591];
                
                r_data[16593] <= r_data[16592];
                
                r_data[16594] <= r_data[16593];
                
                r_data[16595] <= r_data[16594];
                
                r_data[16596] <= r_data[16595];
                
                r_data[16597] <= r_data[16596];
                
                r_data[16598] <= r_data[16597];
                
                r_data[16599] <= r_data[16598];
                
                r_data[16600] <= r_data[16599];
                
                r_data[16601] <= r_data[16600];
                
                r_data[16602] <= r_data[16601];
                
                r_data[16603] <= r_data[16602];
                
                r_data[16604] <= r_data[16603];
                
                r_data[16605] <= r_data[16604];
                
                r_data[16606] <= r_data[16605];
                
                r_data[16607] <= r_data[16606];
                
                r_data[16608] <= r_data[16607];
                
                r_data[16609] <= r_data[16608];
                
                r_data[16610] <= r_data[16609];
                
                r_data[16611] <= r_data[16610];
                
                r_data[16612] <= r_data[16611];
                
                r_data[16613] <= r_data[16612];
                
                r_data[16614] <= r_data[16613];
                
                r_data[16615] <= r_data[16614];
                
                r_data[16616] <= r_data[16615];
                
                r_data[16617] <= r_data[16616];
                
                r_data[16618] <= r_data[16617];
                
                r_data[16619] <= r_data[16618];
                
                r_data[16620] <= r_data[16619];
                
                r_data[16621] <= r_data[16620];
                
                r_data[16622] <= r_data[16621];
                
                r_data[16623] <= r_data[16622];
                
                r_data[16624] <= r_data[16623];
                
                r_data[16625] <= r_data[16624];
                
                r_data[16626] <= r_data[16625];
                
                r_data[16627] <= r_data[16626];
                
                r_data[16628] <= r_data[16627];
                
                r_data[16629] <= r_data[16628];
                
                r_data[16630] <= r_data[16629];
                
                r_data[16631] <= r_data[16630];
                
                r_data[16632] <= r_data[16631];
                
                r_data[16633] <= r_data[16632];
                
                r_data[16634] <= r_data[16633];
                
                r_data[16635] <= r_data[16634];
                
                r_data[16636] <= r_data[16635];
                
                r_data[16637] <= r_data[16636];
                
                r_data[16638] <= r_data[16637];
                
                r_data[16639] <= r_data[16638];
                
                r_data[16640] <= r_data[16639];
                
                r_data[16641] <= r_data[16640];
                
                r_data[16642] <= r_data[16641];
                
                r_data[16643] <= r_data[16642];
                
                r_data[16644] <= r_data[16643];
                
                r_data[16645] <= r_data[16644];
                
                r_data[16646] <= r_data[16645];
                
                r_data[16647] <= r_data[16646];
                
                r_data[16648] <= r_data[16647];
                
                r_data[16649] <= r_data[16648];
                
                r_data[16650] <= r_data[16649];
                
                r_data[16651] <= r_data[16650];
                
                r_data[16652] <= r_data[16651];
                
                r_data[16653] <= r_data[16652];
                
                r_data[16654] <= r_data[16653];
                
                r_data[16655] <= r_data[16654];
                
                r_data[16656] <= r_data[16655];
                
                r_data[16657] <= r_data[16656];
                
                r_data[16658] <= r_data[16657];
                
                r_data[16659] <= r_data[16658];
                
                r_data[16660] <= r_data[16659];
                
                r_data[16661] <= r_data[16660];
                
                r_data[16662] <= r_data[16661];
                
                r_data[16663] <= r_data[16662];
                
                r_data[16664] <= r_data[16663];
                
                r_data[16665] <= r_data[16664];
                
                r_data[16666] <= r_data[16665];
                
                r_data[16667] <= r_data[16666];
                
                r_data[16668] <= r_data[16667];
                
                r_data[16669] <= r_data[16668];
                
                r_data[16670] <= r_data[16669];
                
                r_data[16671] <= r_data[16670];
                
                r_data[16672] <= r_data[16671];
                
                r_data[16673] <= r_data[16672];
                
                r_data[16674] <= r_data[16673];
                
                r_data[16675] <= r_data[16674];
                
                r_data[16676] <= r_data[16675];
                
                r_data[16677] <= r_data[16676];
                
                r_data[16678] <= r_data[16677];
                
                r_data[16679] <= r_data[16678];
                
                r_data[16680] <= r_data[16679];
                
                r_data[16681] <= r_data[16680];
                
                r_data[16682] <= r_data[16681];
                
                r_data[16683] <= r_data[16682];
                
                r_data[16684] <= r_data[16683];
                
                r_data[16685] <= r_data[16684];
                
                r_data[16686] <= r_data[16685];
                
                r_data[16687] <= r_data[16686];
                
                r_data[16688] <= r_data[16687];
                
                r_data[16689] <= r_data[16688];
                
                r_data[16690] <= r_data[16689];
                
                r_data[16691] <= r_data[16690];
                
                r_data[16692] <= r_data[16691];
                
                r_data[16693] <= r_data[16692];
                
                r_data[16694] <= r_data[16693];
                
                r_data[16695] <= r_data[16694];
                
                r_data[16696] <= r_data[16695];
                
                r_data[16697] <= r_data[16696];
                
                r_data[16698] <= r_data[16697];
                
                r_data[16699] <= r_data[16698];
                
                r_data[16700] <= r_data[16699];
                
                r_data[16701] <= r_data[16700];
                
                r_data[16702] <= r_data[16701];
                
                r_data[16703] <= r_data[16702];
                
                r_data[16704] <= r_data[16703];
                
                r_data[16705] <= r_data[16704];
                
                r_data[16706] <= r_data[16705];
                
                r_data[16707] <= r_data[16706];
                
                r_data[16708] <= r_data[16707];
                
                r_data[16709] <= r_data[16708];
                
                r_data[16710] <= r_data[16709];
                
                r_data[16711] <= r_data[16710];
                
                r_data[16712] <= r_data[16711];
                
                r_data[16713] <= r_data[16712];
                
                r_data[16714] <= r_data[16713];
                
                r_data[16715] <= r_data[16714];
                
                r_data[16716] <= r_data[16715];
                
                r_data[16717] <= r_data[16716];
                
                r_data[16718] <= r_data[16717];
                
                r_data[16719] <= r_data[16718];
                
                r_data[16720] <= r_data[16719];
                
                r_data[16721] <= r_data[16720];
                
                r_data[16722] <= r_data[16721];
                
                r_data[16723] <= r_data[16722];
                
                r_data[16724] <= r_data[16723];
                
                r_data[16725] <= r_data[16724];
                
                r_data[16726] <= r_data[16725];
                
                r_data[16727] <= r_data[16726];
                
                r_data[16728] <= r_data[16727];
                
                r_data[16729] <= r_data[16728];
                
                r_data[16730] <= r_data[16729];
                
                r_data[16731] <= r_data[16730];
                
                r_data[16732] <= r_data[16731];
                
                r_data[16733] <= r_data[16732];
                
                r_data[16734] <= r_data[16733];
                
                r_data[16735] <= r_data[16734];
                
                r_data[16736] <= r_data[16735];
                
                r_data[16737] <= r_data[16736];
                
                r_data[16738] <= r_data[16737];
                
                r_data[16739] <= r_data[16738];
                
                r_data[16740] <= r_data[16739];
                
                r_data[16741] <= r_data[16740];
                
                r_data[16742] <= r_data[16741];
                
                r_data[16743] <= r_data[16742];
                
                r_data[16744] <= r_data[16743];
                
                r_data[16745] <= r_data[16744];
                
                r_data[16746] <= r_data[16745];
                
                r_data[16747] <= r_data[16746];
                
                r_data[16748] <= r_data[16747];
                
                r_data[16749] <= r_data[16748];
                
                r_data[16750] <= r_data[16749];
                
                r_data[16751] <= r_data[16750];
                
                r_data[16752] <= r_data[16751];
                
                r_data[16753] <= r_data[16752];
                
                r_data[16754] <= r_data[16753];
                
                r_data[16755] <= r_data[16754];
                
                r_data[16756] <= r_data[16755];
                
                r_data[16757] <= r_data[16756];
                
                r_data[16758] <= r_data[16757];
                
                r_data[16759] <= r_data[16758];
                
                r_data[16760] <= r_data[16759];
                
                r_data[16761] <= r_data[16760];
                
                r_data[16762] <= r_data[16761];
                
                r_data[16763] <= r_data[16762];
                
                r_data[16764] <= r_data[16763];
                
                r_data[16765] <= r_data[16764];
                
                r_data[16766] <= r_data[16765];
                
                r_data[16767] <= r_data[16766];
                
                r_data[16768] <= r_data[16767];
                
                r_data[16769] <= r_data[16768];
                
                r_data[16770] <= r_data[16769];
                
                r_data[16771] <= r_data[16770];
                
                r_data[16772] <= r_data[16771];
                
                r_data[16773] <= r_data[16772];
                
                r_data[16774] <= r_data[16773];
                
                r_data[16775] <= r_data[16774];
                
                r_data[16776] <= r_data[16775];
                
                r_data[16777] <= r_data[16776];
                
                r_data[16778] <= r_data[16777];
                
                r_data[16779] <= r_data[16778];
                
                r_data[16780] <= r_data[16779];
                
                r_data[16781] <= r_data[16780];
                
                r_data[16782] <= r_data[16781];
                
                r_data[16783] <= r_data[16782];
                
                r_data[16784] <= r_data[16783];
                
                r_data[16785] <= r_data[16784];
                
                r_data[16786] <= r_data[16785];
                
                r_data[16787] <= r_data[16786];
                
                r_data[16788] <= r_data[16787];
                
                r_data[16789] <= r_data[16788];
                
                r_data[16790] <= r_data[16789];
                
                r_data[16791] <= r_data[16790];
                
                r_data[16792] <= r_data[16791];
                
                r_data[16793] <= r_data[16792];
                
                r_data[16794] <= r_data[16793];
                
                r_data[16795] <= r_data[16794];
                
                r_data[16796] <= r_data[16795];
                
                r_data[16797] <= r_data[16796];
                
                r_data[16798] <= r_data[16797];
                
                r_data[16799] <= r_data[16798];
                
                r_data[16800] <= r_data[16799];
                
                r_data[16801] <= r_data[16800];
                
                r_data[16802] <= r_data[16801];
                
                r_data[16803] <= r_data[16802];
                
                r_data[16804] <= r_data[16803];
                
                r_data[16805] <= r_data[16804];
                
                r_data[16806] <= r_data[16805];
                
                r_data[16807] <= r_data[16806];
                
                r_data[16808] <= r_data[16807];
                
                r_data[16809] <= r_data[16808];
                
                r_data[16810] <= r_data[16809];
                
                r_data[16811] <= r_data[16810];
                
                r_data[16812] <= r_data[16811];
                
                r_data[16813] <= r_data[16812];
                
                r_data[16814] <= r_data[16813];
                
                r_data[16815] <= r_data[16814];
                
                r_data[16816] <= r_data[16815];
                
                r_data[16817] <= r_data[16816];
                
                r_data[16818] <= r_data[16817];
                
                r_data[16819] <= r_data[16818];
                
                r_data[16820] <= r_data[16819];
                
                r_data[16821] <= r_data[16820];
                
                r_data[16822] <= r_data[16821];
                
                r_data[16823] <= r_data[16822];
                
                r_data[16824] <= r_data[16823];
                
                r_data[16825] <= r_data[16824];
                
                r_data[16826] <= r_data[16825];
                
                r_data[16827] <= r_data[16826];
                
                r_data[16828] <= r_data[16827];
                
                r_data[16829] <= r_data[16828];
                
                r_data[16830] <= r_data[16829];
                
                r_data[16831] <= r_data[16830];
                
                r_data[16832] <= r_data[16831];
                
                r_data[16833] <= r_data[16832];
                
                r_data[16834] <= r_data[16833];
                
                r_data[16835] <= r_data[16834];
                
                r_data[16836] <= r_data[16835];
                
                r_data[16837] <= r_data[16836];
                
                r_data[16838] <= r_data[16837];
                
                r_data[16839] <= r_data[16838];
                
                r_data[16840] <= r_data[16839];
                
                r_data[16841] <= r_data[16840];
                
                r_data[16842] <= r_data[16841];
                
                r_data[16843] <= r_data[16842];
                
                r_data[16844] <= r_data[16843];
                
                r_data[16845] <= r_data[16844];
                
                r_data[16846] <= r_data[16845];
                
                r_data[16847] <= r_data[16846];
                
                r_data[16848] <= r_data[16847];
                
                r_data[16849] <= r_data[16848];
                
                r_data[16850] <= r_data[16849];
                
                r_data[16851] <= r_data[16850];
                
                r_data[16852] <= r_data[16851];
                
                r_data[16853] <= r_data[16852];
                
                r_data[16854] <= r_data[16853];
                
                r_data[16855] <= r_data[16854];
                
                r_data[16856] <= r_data[16855];
                
                r_data[16857] <= r_data[16856];
                
                r_data[16858] <= r_data[16857];
                
                r_data[16859] <= r_data[16858];
                
                r_data[16860] <= r_data[16859];
                
                r_data[16861] <= r_data[16860];
                
                r_data[16862] <= r_data[16861];
                
                r_data[16863] <= r_data[16862];
                
                r_data[16864] <= r_data[16863];
                
                r_data[16865] <= r_data[16864];
                
                r_data[16866] <= r_data[16865];
                
                r_data[16867] <= r_data[16866];
                
                r_data[16868] <= r_data[16867];
                
                r_data[16869] <= r_data[16868];
                
                r_data[16870] <= r_data[16869];
                
                r_data[16871] <= r_data[16870];
                
                r_data[16872] <= r_data[16871];
                
                r_data[16873] <= r_data[16872];
                
                r_data[16874] <= r_data[16873];
                
                r_data[16875] <= r_data[16874];
                
                r_data[16876] <= r_data[16875];
                
                r_data[16877] <= r_data[16876];
                
                r_data[16878] <= r_data[16877];
                
                r_data[16879] <= r_data[16878];
                
                r_data[16880] <= r_data[16879];
                
                r_data[16881] <= r_data[16880];
                
                r_data[16882] <= r_data[16881];
                
                r_data[16883] <= r_data[16882];
                
                r_data[16884] <= r_data[16883];
                
                r_data[16885] <= r_data[16884];
                
                r_data[16886] <= r_data[16885];
                
                r_data[16887] <= r_data[16886];
                
                r_data[16888] <= r_data[16887];
                
                r_data[16889] <= r_data[16888];
                
                r_data[16890] <= r_data[16889];
                
                r_data[16891] <= r_data[16890];
                
                r_data[16892] <= r_data[16891];
                
                r_data[16893] <= r_data[16892];
                
                r_data[16894] <= r_data[16893];
                
                r_data[16895] <= r_data[16894];
                
                r_data[16896] <= r_data[16895];
                
                r_data[16897] <= r_data[16896];
                
                r_data[16898] <= r_data[16897];
                
                r_data[16899] <= r_data[16898];
                
                r_data[16900] <= r_data[16899];
                
                r_data[16901] <= r_data[16900];
                
                r_data[16902] <= r_data[16901];
                
                r_data[16903] <= r_data[16902];
                
                r_data[16904] <= r_data[16903];
                
                r_data[16905] <= r_data[16904];
                
                r_data[16906] <= r_data[16905];
                
                r_data[16907] <= r_data[16906];
                
                r_data[16908] <= r_data[16907];
                
                r_data[16909] <= r_data[16908];
                
                r_data[16910] <= r_data[16909];
                
                r_data[16911] <= r_data[16910];
                
                r_data[16912] <= r_data[16911];
                
                r_data[16913] <= r_data[16912];
                
                r_data[16914] <= r_data[16913];
                
                r_data[16915] <= r_data[16914];
                
                r_data[16916] <= r_data[16915];
                
                r_data[16917] <= r_data[16916];
                
                r_data[16918] <= r_data[16917];
                
                r_data[16919] <= r_data[16918];
                
                r_data[16920] <= r_data[16919];
                
                r_data[16921] <= r_data[16920];
                
                r_data[16922] <= r_data[16921];
                
                r_data[16923] <= r_data[16922];
                
                r_data[16924] <= r_data[16923];
                
                r_data[16925] <= r_data[16924];
                
                r_data[16926] <= r_data[16925];
                
                r_data[16927] <= r_data[16926];
                
                r_data[16928] <= r_data[16927];
                
                r_data[16929] <= r_data[16928];
                
                r_data[16930] <= r_data[16929];
                
                r_data[16931] <= r_data[16930];
                
                r_data[16932] <= r_data[16931];
                
                r_data[16933] <= r_data[16932];
                
                r_data[16934] <= r_data[16933];
                
                r_data[16935] <= r_data[16934];
                
                r_data[16936] <= r_data[16935];
                
                r_data[16937] <= r_data[16936];
                
                r_data[16938] <= r_data[16937];
                
                r_data[16939] <= r_data[16938];
                
                r_data[16940] <= r_data[16939];
                
                r_data[16941] <= r_data[16940];
                
                r_data[16942] <= r_data[16941];
                
                r_data[16943] <= r_data[16942];
                
                r_data[16944] <= r_data[16943];
                
                r_data[16945] <= r_data[16944];
                
                r_data[16946] <= r_data[16945];
                
                r_data[16947] <= r_data[16946];
                
                r_data[16948] <= r_data[16947];
                
                r_data[16949] <= r_data[16948];
                
                r_data[16950] <= r_data[16949];
                
                r_data[16951] <= r_data[16950];
                
                r_data[16952] <= r_data[16951];
                
                r_data[16953] <= r_data[16952];
                
                r_data[16954] <= r_data[16953];
                
                r_data[16955] <= r_data[16954];
                
                r_data[16956] <= r_data[16955];
                
                r_data[16957] <= r_data[16956];
                
                r_data[16958] <= r_data[16957];
                
                r_data[16959] <= r_data[16958];
                
                r_data[16960] <= r_data[16959];
                
                r_data[16961] <= r_data[16960];
                
                r_data[16962] <= r_data[16961];
                
                r_data[16963] <= r_data[16962];
                
                r_data[16964] <= r_data[16963];
                
                r_data[16965] <= r_data[16964];
                
                r_data[16966] <= r_data[16965];
                
                r_data[16967] <= r_data[16966];
                
                r_data[16968] <= r_data[16967];
                
                r_data[16969] <= r_data[16968];
                
                r_data[16970] <= r_data[16969];
                
                r_data[16971] <= r_data[16970];
                
                r_data[16972] <= r_data[16971];
                
                r_data[16973] <= r_data[16972];
                
                r_data[16974] <= r_data[16973];
                
                r_data[16975] <= r_data[16974];
                
                r_data[16976] <= r_data[16975];
                
                r_data[16977] <= r_data[16976];
                
                r_data[16978] <= r_data[16977];
                
                r_data[16979] <= r_data[16978];
                
                r_data[16980] <= r_data[16979];
                
                r_data[16981] <= r_data[16980];
                
                r_data[16982] <= r_data[16981];
                
                r_data[16983] <= r_data[16982];
                
                r_data[16984] <= r_data[16983];
                
                r_data[16985] <= r_data[16984];
                
                r_data[16986] <= r_data[16985];
                
                r_data[16987] <= r_data[16986];
                
                r_data[16988] <= r_data[16987];
                
                r_data[16989] <= r_data[16988];
                
                r_data[16990] <= r_data[16989];
                
                r_data[16991] <= r_data[16990];
                
                r_data[16992] <= r_data[16991];
                
                r_data[16993] <= r_data[16992];
                
                r_data[16994] <= r_data[16993];
                
                r_data[16995] <= r_data[16994];
                
                r_data[16996] <= r_data[16995];
                
                r_data[16997] <= r_data[16996];
                
                r_data[16998] <= r_data[16997];
                
                r_data[16999] <= r_data[16998];
                
                r_data[17000] <= r_data[16999];
                
                r_data[17001] <= r_data[17000];
                
                r_data[17002] <= r_data[17001];
                
                r_data[17003] <= r_data[17002];
                
                r_data[17004] <= r_data[17003];
                
                r_data[17005] <= r_data[17004];
                
                r_data[17006] <= r_data[17005];
                
                r_data[17007] <= r_data[17006];
                
                r_data[17008] <= r_data[17007];
                
                r_data[17009] <= r_data[17008];
                
                r_data[17010] <= r_data[17009];
                
                r_data[17011] <= r_data[17010];
                
                r_data[17012] <= r_data[17011];
                
                r_data[17013] <= r_data[17012];
                
                r_data[17014] <= r_data[17013];
                
                r_data[17015] <= r_data[17014];
                
                r_data[17016] <= r_data[17015];
                
                r_data[17017] <= r_data[17016];
                
                r_data[17018] <= r_data[17017];
                
                r_data[17019] <= r_data[17018];
                
                r_data[17020] <= r_data[17019];
                
                r_data[17021] <= r_data[17020];
                
                r_data[17022] <= r_data[17021];
                
                r_data[17023] <= r_data[17022];
                
                r_data[17024] <= r_data[17023];
                
                r_data[17025] <= r_data[17024];
                
                r_data[17026] <= r_data[17025];
                
                r_data[17027] <= r_data[17026];
                
                r_data[17028] <= r_data[17027];
                
                r_data[17029] <= r_data[17028];
                
                r_data[17030] <= r_data[17029];
                
                r_data[17031] <= r_data[17030];
                
                r_data[17032] <= r_data[17031];
                
                r_data[17033] <= r_data[17032];
                
                r_data[17034] <= r_data[17033];
                
                r_data[17035] <= r_data[17034];
                
                r_data[17036] <= r_data[17035];
                
                r_data[17037] <= r_data[17036];
                
                r_data[17038] <= r_data[17037];
                
                r_data[17039] <= r_data[17038];
                
                r_data[17040] <= r_data[17039];
                
                r_data[17041] <= r_data[17040];
                
                r_data[17042] <= r_data[17041];
                
                r_data[17043] <= r_data[17042];
                
                r_data[17044] <= r_data[17043];
                
                r_data[17045] <= r_data[17044];
                
                r_data[17046] <= r_data[17045];
                
                r_data[17047] <= r_data[17046];
                
                r_data[17048] <= r_data[17047];
                
                r_data[17049] <= r_data[17048];
                
                r_data[17050] <= r_data[17049];
                
                r_data[17051] <= r_data[17050];
                
                r_data[17052] <= r_data[17051];
                
                r_data[17053] <= r_data[17052];
                
                r_data[17054] <= r_data[17053];
                
                r_data[17055] <= r_data[17054];
                
                r_data[17056] <= r_data[17055];
                
                r_data[17057] <= r_data[17056];
                
                r_data[17058] <= r_data[17057];
                
                r_data[17059] <= r_data[17058];
                
                r_data[17060] <= r_data[17059];
                
                r_data[17061] <= r_data[17060];
                
                r_data[17062] <= r_data[17061];
                
                r_data[17063] <= r_data[17062];
                
                r_data[17064] <= r_data[17063];
                
                r_data[17065] <= r_data[17064];
                
                r_data[17066] <= r_data[17065];
                
                r_data[17067] <= r_data[17066];
                
                r_data[17068] <= r_data[17067];
                
                r_data[17069] <= r_data[17068];
                
                r_data[17070] <= r_data[17069];
                
                r_data[17071] <= r_data[17070];
                
                r_data[17072] <= r_data[17071];
                
                r_data[17073] <= r_data[17072];
                
                r_data[17074] <= r_data[17073];
                
                r_data[17075] <= r_data[17074];
                
                r_data[17076] <= r_data[17075];
                
                r_data[17077] <= r_data[17076];
                
                r_data[17078] <= r_data[17077];
                
                r_data[17079] <= r_data[17078];
                
                r_data[17080] <= r_data[17079];
                
                r_data[17081] <= r_data[17080];
                
                r_data[17082] <= r_data[17081];
                
                r_data[17083] <= r_data[17082];
                
                r_data[17084] <= r_data[17083];
                
                r_data[17085] <= r_data[17084];
                
                r_data[17086] <= r_data[17085];
                
                r_data[17087] <= r_data[17086];
                
                r_data[17088] <= r_data[17087];
                
                r_data[17089] <= r_data[17088];
                
                r_data[17090] <= r_data[17089];
                
                r_data[17091] <= r_data[17090];
                
                r_data[17092] <= r_data[17091];
                
                r_data[17093] <= r_data[17092];
                
                r_data[17094] <= r_data[17093];
                
                r_data[17095] <= r_data[17094];
                
                r_data[17096] <= r_data[17095];
                
                r_data[17097] <= r_data[17096];
                
                r_data[17098] <= r_data[17097];
                
                r_data[17099] <= r_data[17098];
                
                r_data[17100] <= r_data[17099];
                
                r_data[17101] <= r_data[17100];
                
                r_data[17102] <= r_data[17101];
                
                r_data[17103] <= r_data[17102];
                
                r_data[17104] <= r_data[17103];
                
                r_data[17105] <= r_data[17104];
                
                r_data[17106] <= r_data[17105];
                
                r_data[17107] <= r_data[17106];
                
                r_data[17108] <= r_data[17107];
                
                r_data[17109] <= r_data[17108];
                
                r_data[17110] <= r_data[17109];
                
                r_data[17111] <= r_data[17110];
                
                r_data[17112] <= r_data[17111];
                
                r_data[17113] <= r_data[17112];
                
                r_data[17114] <= r_data[17113];
                
                r_data[17115] <= r_data[17114];
                
                r_data[17116] <= r_data[17115];
                
                r_data[17117] <= r_data[17116];
                
                r_data[17118] <= r_data[17117];
                
                r_data[17119] <= r_data[17118];
                
                r_data[17120] <= r_data[17119];
                
                r_data[17121] <= r_data[17120];
                
                r_data[17122] <= r_data[17121];
                
                r_data[17123] <= r_data[17122];
                
                r_data[17124] <= r_data[17123];
                
                r_data[17125] <= r_data[17124];
                
                r_data[17126] <= r_data[17125];
                
                r_data[17127] <= r_data[17126];
                
                r_data[17128] <= r_data[17127];
                
                r_data[17129] <= r_data[17128];
                
                r_data[17130] <= r_data[17129];
                
                r_data[17131] <= r_data[17130];
                
                r_data[17132] <= r_data[17131];
                
                r_data[17133] <= r_data[17132];
                
                r_data[17134] <= r_data[17133];
                
                r_data[17135] <= r_data[17134];
                
                r_data[17136] <= r_data[17135];
                
                r_data[17137] <= r_data[17136];
                
                r_data[17138] <= r_data[17137];
                
                r_data[17139] <= r_data[17138];
                
                r_data[17140] <= r_data[17139];
                
                r_data[17141] <= r_data[17140];
                
                r_data[17142] <= r_data[17141];
                
                r_data[17143] <= r_data[17142];
                
                r_data[17144] <= r_data[17143];
                
                r_data[17145] <= r_data[17144];
                
                r_data[17146] <= r_data[17145];
                
                r_data[17147] <= r_data[17146];
                
                r_data[17148] <= r_data[17147];
                
                r_data[17149] <= r_data[17148];
                
                r_data[17150] <= r_data[17149];
                
                r_data[17151] <= r_data[17150];
                
                r_data[17152] <= r_data[17151];
                
                r_data[17153] <= r_data[17152];
                
                r_data[17154] <= r_data[17153];
                
                r_data[17155] <= r_data[17154];
                
                r_data[17156] <= r_data[17155];
                
                r_data[17157] <= r_data[17156];
                
                r_data[17158] <= r_data[17157];
                
                r_data[17159] <= r_data[17158];
                
                r_data[17160] <= r_data[17159];
                
                r_data[17161] <= r_data[17160];
                
                r_data[17162] <= r_data[17161];
                
                r_data[17163] <= r_data[17162];
                
                r_data[17164] <= r_data[17163];
                
                r_data[17165] <= r_data[17164];
                
                r_data[17166] <= r_data[17165];
                
                r_data[17167] <= r_data[17166];
                
                r_data[17168] <= r_data[17167];
                
                r_data[17169] <= r_data[17168];
                
                r_data[17170] <= r_data[17169];
                
                r_data[17171] <= r_data[17170];
                
                r_data[17172] <= r_data[17171];
                
                r_data[17173] <= r_data[17172];
                
                r_data[17174] <= r_data[17173];
                
                r_data[17175] <= r_data[17174];
                
                r_data[17176] <= r_data[17175];
                
                r_data[17177] <= r_data[17176];
                
                r_data[17178] <= r_data[17177];
                
                r_data[17179] <= r_data[17178];
                
                r_data[17180] <= r_data[17179];
                
                r_data[17181] <= r_data[17180];
                
                r_data[17182] <= r_data[17181];
                
                r_data[17183] <= r_data[17182];
                
                r_data[17184] <= r_data[17183];
                
                r_data[17185] <= r_data[17184];
                
                r_data[17186] <= r_data[17185];
                
                r_data[17187] <= r_data[17186];
                
                r_data[17188] <= r_data[17187];
                
                r_data[17189] <= r_data[17188];
                
                r_data[17190] <= r_data[17189];
                
                r_data[17191] <= r_data[17190];
                
                r_data[17192] <= r_data[17191];
                
                r_data[17193] <= r_data[17192];
                
                r_data[17194] <= r_data[17193];
                
                r_data[17195] <= r_data[17194];
                
                r_data[17196] <= r_data[17195];
                
                r_data[17197] <= r_data[17196];
                
                r_data[17198] <= r_data[17197];
                
                r_data[17199] <= r_data[17198];
                
                r_data[17200] <= r_data[17199];
                
                r_data[17201] <= r_data[17200];
                
                r_data[17202] <= r_data[17201];
                
                r_data[17203] <= r_data[17202];
                
                r_data[17204] <= r_data[17203];
                
                r_data[17205] <= r_data[17204];
                
                r_data[17206] <= r_data[17205];
                
                r_data[17207] <= r_data[17206];
                
                r_data[17208] <= r_data[17207];
                
                r_data[17209] <= r_data[17208];
                
                r_data[17210] <= r_data[17209];
                
                r_data[17211] <= r_data[17210];
                
                r_data[17212] <= r_data[17211];
                
                r_data[17213] <= r_data[17212];
                
                r_data[17214] <= r_data[17213];
                
                r_data[17215] <= r_data[17214];
                
                r_data[17216] <= r_data[17215];
                
                r_data[17217] <= r_data[17216];
                
                r_data[17218] <= r_data[17217];
                
                r_data[17219] <= r_data[17218];
                
                r_data[17220] <= r_data[17219];
                
                r_data[17221] <= r_data[17220];
                
                r_data[17222] <= r_data[17221];
                
                r_data[17223] <= r_data[17222];
                
                r_data[17224] <= r_data[17223];
                
                r_data[17225] <= r_data[17224];
                
                r_data[17226] <= r_data[17225];
                
                r_data[17227] <= r_data[17226];
                
                r_data[17228] <= r_data[17227];
                
                r_data[17229] <= r_data[17228];
                
                r_data[17230] <= r_data[17229];
                
                r_data[17231] <= r_data[17230];
                
                r_data[17232] <= r_data[17231];
                
                r_data[17233] <= r_data[17232];
                
                r_data[17234] <= r_data[17233];
                
                r_data[17235] <= r_data[17234];
                
                r_data[17236] <= r_data[17235];
                
                r_data[17237] <= r_data[17236];
                
                r_data[17238] <= r_data[17237];
                
                r_data[17239] <= r_data[17238];
                
                r_data[17240] <= r_data[17239];
                
                r_data[17241] <= r_data[17240];
                
                r_data[17242] <= r_data[17241];
                
                r_data[17243] <= r_data[17242];
                
                r_data[17244] <= r_data[17243];
                
                r_data[17245] <= r_data[17244];
                
                r_data[17246] <= r_data[17245];
                
                r_data[17247] <= r_data[17246];
                
                r_data[17248] <= r_data[17247];
                
                r_data[17249] <= r_data[17248];
                
                r_data[17250] <= r_data[17249];
                
                r_data[17251] <= r_data[17250];
                
                r_data[17252] <= r_data[17251];
                
                r_data[17253] <= r_data[17252];
                
                r_data[17254] <= r_data[17253];
                
                r_data[17255] <= r_data[17254];
                
                r_data[17256] <= r_data[17255];
                
                r_data[17257] <= r_data[17256];
                
                r_data[17258] <= r_data[17257];
                
                r_data[17259] <= r_data[17258];
                
                r_data[17260] <= r_data[17259];
                
                r_data[17261] <= r_data[17260];
                
                r_data[17262] <= r_data[17261];
                
                r_data[17263] <= r_data[17262];
                
                r_data[17264] <= r_data[17263];
                
                r_data[17265] <= r_data[17264];
                
                r_data[17266] <= r_data[17265];
                
                r_data[17267] <= r_data[17266];
                
                r_data[17268] <= r_data[17267];
                
                r_data[17269] <= r_data[17268];
                
                r_data[17270] <= r_data[17269];
                
                r_data[17271] <= r_data[17270];
                
                r_data[17272] <= r_data[17271];
                
                r_data[17273] <= r_data[17272];
                
                r_data[17274] <= r_data[17273];
                
                r_data[17275] <= r_data[17274];
                
                r_data[17276] <= r_data[17275];
                
                r_data[17277] <= r_data[17276];
                
                r_data[17278] <= r_data[17277];
                
                r_data[17279] <= r_data[17278];
                
                r_data[17280] <= r_data[17279];
                
                r_data[17281] <= r_data[17280];
                
                r_data[17282] <= r_data[17281];
                
                r_data[17283] <= r_data[17282];
                
                r_data[17284] <= r_data[17283];
                
                r_data[17285] <= r_data[17284];
                
                r_data[17286] <= r_data[17285];
                
                r_data[17287] <= r_data[17286];
                
                r_data[17288] <= r_data[17287];
                
                r_data[17289] <= r_data[17288];
                
                r_data[17290] <= r_data[17289];
                
                r_data[17291] <= r_data[17290];
                
                r_data[17292] <= r_data[17291];
                
                r_data[17293] <= r_data[17292];
                
                r_data[17294] <= r_data[17293];
                
                r_data[17295] <= r_data[17294];
                
                r_data[17296] <= r_data[17295];
                
                r_data[17297] <= r_data[17296];
                
                r_data[17298] <= r_data[17297];
                
                r_data[17299] <= r_data[17298];
                
                r_data[17300] <= r_data[17299];
                
                r_data[17301] <= r_data[17300];
                
                r_data[17302] <= r_data[17301];
                
                r_data[17303] <= r_data[17302];
                
                r_data[17304] <= r_data[17303];
                
                r_data[17305] <= r_data[17304];
                
                r_data[17306] <= r_data[17305];
                
                r_data[17307] <= r_data[17306];
                
                r_data[17308] <= r_data[17307];
                
                r_data[17309] <= r_data[17308];
                
                r_data[17310] <= r_data[17309];
                
                r_data[17311] <= r_data[17310];
                
                r_data[17312] <= r_data[17311];
                
                r_data[17313] <= r_data[17312];
                
                r_data[17314] <= r_data[17313];
                
                r_data[17315] <= r_data[17314];
                
                r_data[17316] <= r_data[17315];
                
                r_data[17317] <= r_data[17316];
                
                r_data[17318] <= r_data[17317];
                
                r_data[17319] <= r_data[17318];
                
                r_data[17320] <= r_data[17319];
                
                r_data[17321] <= r_data[17320];
                
                r_data[17322] <= r_data[17321];
                
                r_data[17323] <= r_data[17322];
                
                r_data[17324] <= r_data[17323];
                
                r_data[17325] <= r_data[17324];
                
                r_data[17326] <= r_data[17325];
                
                r_data[17327] <= r_data[17326];
                
                r_data[17328] <= r_data[17327];
                
                r_data[17329] <= r_data[17328];
                
                r_data[17330] <= r_data[17329];
                
                r_data[17331] <= r_data[17330];
                
                r_data[17332] <= r_data[17331];
                
                r_data[17333] <= r_data[17332];
                
                r_data[17334] <= r_data[17333];
                
                r_data[17335] <= r_data[17334];
                
                r_data[17336] <= r_data[17335];
                
                r_data[17337] <= r_data[17336];
                
                r_data[17338] <= r_data[17337];
                
                r_data[17339] <= r_data[17338];
                
                r_data[17340] <= r_data[17339];
                
                r_data[17341] <= r_data[17340];
                
                r_data[17342] <= r_data[17341];
                
                r_data[17343] <= r_data[17342];
                
                r_data[17344] <= r_data[17343];
                
                r_data[17345] <= r_data[17344];
                
                r_data[17346] <= r_data[17345];
                
                r_data[17347] <= r_data[17346];
                
                r_data[17348] <= r_data[17347];
                
                r_data[17349] <= r_data[17348];
                
                r_data[17350] <= r_data[17349];
                
                r_data[17351] <= r_data[17350];
                
                r_data[17352] <= r_data[17351];
                
                r_data[17353] <= r_data[17352];
                
                r_data[17354] <= r_data[17353];
                
                r_data[17355] <= r_data[17354];
                
                r_data[17356] <= r_data[17355];
                
                r_data[17357] <= r_data[17356];
                
                r_data[17358] <= r_data[17357];
                
                r_data[17359] <= r_data[17358];
                
                r_data[17360] <= r_data[17359];
                
                r_data[17361] <= r_data[17360];
                
                r_data[17362] <= r_data[17361];
                
                r_data[17363] <= r_data[17362];
                
                r_data[17364] <= r_data[17363];
                
                r_data[17365] <= r_data[17364];
                
                r_data[17366] <= r_data[17365];
                
                r_data[17367] <= r_data[17366];
                
                r_data[17368] <= r_data[17367];
                
                r_data[17369] <= r_data[17368];
                
                r_data[17370] <= r_data[17369];
                
                r_data[17371] <= r_data[17370];
                
                r_data[17372] <= r_data[17371];
                
                r_data[17373] <= r_data[17372];
                
                r_data[17374] <= r_data[17373];
                
                r_data[17375] <= r_data[17374];
                
                r_data[17376] <= r_data[17375];
                
                r_data[17377] <= r_data[17376];
                
                r_data[17378] <= r_data[17377];
                
                r_data[17379] <= r_data[17378];
                
                r_data[17380] <= r_data[17379];
                
                r_data[17381] <= r_data[17380];
                
                r_data[17382] <= r_data[17381];
                
                r_data[17383] <= r_data[17382];
                
                r_data[17384] <= r_data[17383];
                
                r_data[17385] <= r_data[17384];
                
                r_data[17386] <= r_data[17385];
                
                r_data[17387] <= r_data[17386];
                
                r_data[17388] <= r_data[17387];
                
                r_data[17389] <= r_data[17388];
                
                r_data[17390] <= r_data[17389];
                
                r_data[17391] <= r_data[17390];
                
                r_data[17392] <= r_data[17391];
                
                r_data[17393] <= r_data[17392];
                
                r_data[17394] <= r_data[17393];
                
                r_data[17395] <= r_data[17394];
                
                r_data[17396] <= r_data[17395];
                
                r_data[17397] <= r_data[17396];
                
                r_data[17398] <= r_data[17397];
                
                r_data[17399] <= r_data[17398];
                
                r_data[17400] <= r_data[17399];
                
                r_data[17401] <= r_data[17400];
                
                r_data[17402] <= r_data[17401];
                
                r_data[17403] <= r_data[17402];
                
                r_data[17404] <= r_data[17403];
                
                r_data[17405] <= r_data[17404];
                
                r_data[17406] <= r_data[17405];
                
                r_data[17407] <= r_data[17406];
                
                r_data[17408] <= r_data[17407];
                
                r_data[17409] <= r_data[17408];
                
                r_data[17410] <= r_data[17409];
                
                r_data[17411] <= r_data[17410];
                
                r_data[17412] <= r_data[17411];
                
                r_data[17413] <= r_data[17412];
                
                r_data[17414] <= r_data[17413];
                
                r_data[17415] <= r_data[17414];
                
                r_data[17416] <= r_data[17415];
                
                r_data[17417] <= r_data[17416];
                
                r_data[17418] <= r_data[17417];
                
                r_data[17419] <= r_data[17418];
                
                r_data[17420] <= r_data[17419];
                
                r_data[17421] <= r_data[17420];
                
                r_data[17422] <= r_data[17421];
                
                r_data[17423] <= r_data[17422];
                
                r_data[17424] <= r_data[17423];
                
                r_data[17425] <= r_data[17424];
                
                r_data[17426] <= r_data[17425];
                
                r_data[17427] <= r_data[17426];
                
                r_data[17428] <= r_data[17427];
                
                r_data[17429] <= r_data[17428];
                
                r_data[17430] <= r_data[17429];
                
                r_data[17431] <= r_data[17430];
                
                r_data[17432] <= r_data[17431];
                
                r_data[17433] <= r_data[17432];
                
                r_data[17434] <= r_data[17433];
                
                r_data[17435] <= r_data[17434];
                
                r_data[17436] <= r_data[17435];
                
                r_data[17437] <= r_data[17436];
                
                r_data[17438] <= r_data[17437];
                
                r_data[17439] <= r_data[17438];
                
                r_data[17440] <= r_data[17439];
                
                r_data[17441] <= r_data[17440];
                
                r_data[17442] <= r_data[17441];
                
                r_data[17443] <= r_data[17442];
                
                r_data[17444] <= r_data[17443];
                
                r_data[17445] <= r_data[17444];
                
                r_data[17446] <= r_data[17445];
                
                r_data[17447] <= r_data[17446];
                
                r_data[17448] <= r_data[17447];
                
                r_data[17449] <= r_data[17448];
                
                r_data[17450] <= r_data[17449];
                
                r_data[17451] <= r_data[17450];
                
                r_data[17452] <= r_data[17451];
                
                r_data[17453] <= r_data[17452];
                
                r_data[17454] <= r_data[17453];
                
                r_data[17455] <= r_data[17454];
                
                r_data[17456] <= r_data[17455];
                
                r_data[17457] <= r_data[17456];
                
                r_data[17458] <= r_data[17457];
                
                r_data[17459] <= r_data[17458];
                
                r_data[17460] <= r_data[17459];
                
                r_data[17461] <= r_data[17460];
                
                r_data[17462] <= r_data[17461];
                
                r_data[17463] <= r_data[17462];
                
                r_data[17464] <= r_data[17463];
                
                r_data[17465] <= r_data[17464];
                
                r_data[17466] <= r_data[17465];
                
                r_data[17467] <= r_data[17466];
                
                r_data[17468] <= r_data[17467];
                
                r_data[17469] <= r_data[17468];
                
                r_data[17470] <= r_data[17469];
                
                r_data[17471] <= r_data[17470];
                
                r_data[17472] <= r_data[17471];
                
                r_data[17473] <= r_data[17472];
                
                r_data[17474] <= r_data[17473];
                
                r_data[17475] <= r_data[17474];
                
                r_data[17476] <= r_data[17475];
                
                r_data[17477] <= r_data[17476];
                
                r_data[17478] <= r_data[17477];
                
                r_data[17479] <= r_data[17478];
                
                r_data[17480] <= r_data[17479];
                
                r_data[17481] <= r_data[17480];
                
                r_data[17482] <= r_data[17481];
                
                r_data[17483] <= r_data[17482];
                
                r_data[17484] <= r_data[17483];
                
                r_data[17485] <= r_data[17484];
                
                r_data[17486] <= r_data[17485];
                
                r_data[17487] <= r_data[17486];
                
                r_data[17488] <= r_data[17487];
                
                r_data[17489] <= r_data[17488];
                
                r_data[17490] <= r_data[17489];
                
                r_data[17491] <= r_data[17490];
                
                r_data[17492] <= r_data[17491];
                
                r_data[17493] <= r_data[17492];
                
                r_data[17494] <= r_data[17493];
                
                r_data[17495] <= r_data[17494];
                
                r_data[17496] <= r_data[17495];
                
                r_data[17497] <= r_data[17496];
                
                r_data[17498] <= r_data[17497];
                
                r_data[17499] <= r_data[17498];
                
                r_data[17500] <= r_data[17499];
                
                r_data[17501] <= r_data[17500];
                
                r_data[17502] <= r_data[17501];
                
                r_data[17503] <= r_data[17502];
                
                r_data[17504] <= r_data[17503];
                
                r_data[17505] <= r_data[17504];
                
                r_data[17506] <= r_data[17505];
                
                r_data[17507] <= r_data[17506];
                
                r_data[17508] <= r_data[17507];
                
                r_data[17509] <= r_data[17508];
                
                r_data[17510] <= r_data[17509];
                
                r_data[17511] <= r_data[17510];
                
                r_data[17512] <= r_data[17511];
                
                r_data[17513] <= r_data[17512];
                
                r_data[17514] <= r_data[17513];
                
                r_data[17515] <= r_data[17514];
                
                r_data[17516] <= r_data[17515];
                
                r_data[17517] <= r_data[17516];
                
                r_data[17518] <= r_data[17517];
                
                r_data[17519] <= r_data[17518];
                
                r_data[17520] <= r_data[17519];
                
                r_data[17521] <= r_data[17520];
                
                r_data[17522] <= r_data[17521];
                
                r_data[17523] <= r_data[17522];
                
                r_data[17524] <= r_data[17523];
                
                r_data[17525] <= r_data[17524];
                
                r_data[17526] <= r_data[17525];
                
                r_data[17527] <= r_data[17526];
                
                r_data[17528] <= r_data[17527];
                
                r_data[17529] <= r_data[17528];
                
                r_data[17530] <= r_data[17529];
                
                r_data[17531] <= r_data[17530];
                
                r_data[17532] <= r_data[17531];
                
                r_data[17533] <= r_data[17532];
                
                r_data[17534] <= r_data[17533];
                
                r_data[17535] <= r_data[17534];
                
                r_data[17536] <= r_data[17535];
                
                r_data[17537] <= r_data[17536];
                
                r_data[17538] <= r_data[17537];
                
                r_data[17539] <= r_data[17538];
                
                r_data[17540] <= r_data[17539];
                
                r_data[17541] <= r_data[17540];
                
                r_data[17542] <= r_data[17541];
                
                r_data[17543] <= r_data[17542];
                
                r_data[17544] <= r_data[17543];
                
                r_data[17545] <= r_data[17544];
                
                r_data[17546] <= r_data[17545];
                
                r_data[17547] <= r_data[17546];
                
                r_data[17548] <= r_data[17547];
                
                r_data[17549] <= r_data[17548];
                
                r_data[17550] <= r_data[17549];
                
                r_data[17551] <= r_data[17550];
                
                r_data[17552] <= r_data[17551];
                
                r_data[17553] <= r_data[17552];
                
                r_data[17554] <= r_data[17553];
                
                r_data[17555] <= r_data[17554];
                
                r_data[17556] <= r_data[17555];
                
                r_data[17557] <= r_data[17556];
                
                r_data[17558] <= r_data[17557];
                
                r_data[17559] <= r_data[17558];
                
                r_data[17560] <= r_data[17559];
                
                r_data[17561] <= r_data[17560];
                
                r_data[17562] <= r_data[17561];
                
                r_data[17563] <= r_data[17562];
                
                r_data[17564] <= r_data[17563];
                
                r_data[17565] <= r_data[17564];
                
                r_data[17566] <= r_data[17565];
                
                r_data[17567] <= r_data[17566];
                
                r_data[17568] <= r_data[17567];
                
                r_data[17569] <= r_data[17568];
                
                r_data[17570] <= r_data[17569];
                
                r_data[17571] <= r_data[17570];
                
                r_data[17572] <= r_data[17571];
                
                r_data[17573] <= r_data[17572];
                
                r_data[17574] <= r_data[17573];
                
                r_data[17575] <= r_data[17574];
                
                r_data[17576] <= r_data[17575];
                
                r_data[17577] <= r_data[17576];
                
                r_data[17578] <= r_data[17577];
                
                r_data[17579] <= r_data[17578];
                
                r_data[17580] <= r_data[17579];
                
                r_data[17581] <= r_data[17580];
                
                r_data[17582] <= r_data[17581];
                
                r_data[17583] <= r_data[17582];
                
                r_data[17584] <= r_data[17583];
                
                r_data[17585] <= r_data[17584];
                
                r_data[17586] <= r_data[17585];
                
                r_data[17587] <= r_data[17586];
                
                r_data[17588] <= r_data[17587];
                
                r_data[17589] <= r_data[17588];
                
                r_data[17590] <= r_data[17589];
                
                r_data[17591] <= r_data[17590];
                
                r_data[17592] <= r_data[17591];
                
                r_data[17593] <= r_data[17592];
                
                r_data[17594] <= r_data[17593];
                
                r_data[17595] <= r_data[17594];
                
                r_data[17596] <= r_data[17595];
                
                r_data[17597] <= r_data[17596];
                
                r_data[17598] <= r_data[17597];
                
                r_data[17599] <= r_data[17598];
                
                r_data[17600] <= r_data[17599];
                
                r_data[17601] <= r_data[17600];
                
                r_data[17602] <= r_data[17601];
                
                r_data[17603] <= r_data[17602];
                
                r_data[17604] <= r_data[17603];
                
                r_data[17605] <= r_data[17604];
                
                r_data[17606] <= r_data[17605];
                
                r_data[17607] <= r_data[17606];
                
                r_data[17608] <= r_data[17607];
                
                r_data[17609] <= r_data[17608];
                
                r_data[17610] <= r_data[17609];
                
                r_data[17611] <= r_data[17610];
                
                r_data[17612] <= r_data[17611];
                
                r_data[17613] <= r_data[17612];
                
                r_data[17614] <= r_data[17613];
                
                r_data[17615] <= r_data[17614];
                
                r_data[17616] <= r_data[17615];
                
                r_data[17617] <= r_data[17616];
                
                r_data[17618] <= r_data[17617];
                
                r_data[17619] <= r_data[17618];
                
                r_data[17620] <= r_data[17619];
                
                r_data[17621] <= r_data[17620];
                
                r_data[17622] <= r_data[17621];
                
                r_data[17623] <= r_data[17622];
                
                r_data[17624] <= r_data[17623];
                
                r_data[17625] <= r_data[17624];
                
                r_data[17626] <= r_data[17625];
                
                r_data[17627] <= r_data[17626];
                
                r_data[17628] <= r_data[17627];
                
                r_data[17629] <= r_data[17628];
                
                r_data[17630] <= r_data[17629];
                
                r_data[17631] <= r_data[17630];
                
                r_data[17632] <= r_data[17631];
                
                r_data[17633] <= r_data[17632];
                
                r_data[17634] <= r_data[17633];
                
                r_data[17635] <= r_data[17634];
                
                r_data[17636] <= r_data[17635];
                
                r_data[17637] <= r_data[17636];
                
                r_data[17638] <= r_data[17637];
                
                r_data[17639] <= r_data[17638];
                
                r_data[17640] <= r_data[17639];
                
                r_data[17641] <= r_data[17640];
                
                r_data[17642] <= r_data[17641];
                
                r_data[17643] <= r_data[17642];
                
                r_data[17644] <= r_data[17643];
                
                r_data[17645] <= r_data[17644];
                
                r_data[17646] <= r_data[17645];
                
                r_data[17647] <= r_data[17646];
                
                r_data[17648] <= r_data[17647];
                
                r_data[17649] <= r_data[17648];
                
                r_data[17650] <= r_data[17649];
                
                r_data[17651] <= r_data[17650];
                
                r_data[17652] <= r_data[17651];
                
                r_data[17653] <= r_data[17652];
                
                r_data[17654] <= r_data[17653];
                
                r_data[17655] <= r_data[17654];
                
                r_data[17656] <= r_data[17655];
                
                r_data[17657] <= r_data[17656];
                
                r_data[17658] <= r_data[17657];
                
                r_data[17659] <= r_data[17658];
                
                r_data[17660] <= r_data[17659];
                
                r_data[17661] <= r_data[17660];
                
                r_data[17662] <= r_data[17661];
                
                r_data[17663] <= r_data[17662];
                
                r_data[17664] <= r_data[17663];
                
                r_data[17665] <= r_data[17664];
                
                r_data[17666] <= r_data[17665];
                
                r_data[17667] <= r_data[17666];
                
                r_data[17668] <= r_data[17667];
                
                r_data[17669] <= r_data[17668];
                
                r_data[17670] <= r_data[17669];
                
                r_data[17671] <= r_data[17670];
                
                r_data[17672] <= r_data[17671];
                
                r_data[17673] <= r_data[17672];
                
                r_data[17674] <= r_data[17673];
                
                r_data[17675] <= r_data[17674];
                
                r_data[17676] <= r_data[17675];
                
                r_data[17677] <= r_data[17676];
                
                r_data[17678] <= r_data[17677];
                
                r_data[17679] <= r_data[17678];
                
                r_data[17680] <= r_data[17679];
                
                r_data[17681] <= r_data[17680];
                
                r_data[17682] <= r_data[17681];
                
                r_data[17683] <= r_data[17682];
                
                r_data[17684] <= r_data[17683];
                
                r_data[17685] <= r_data[17684];
                
                r_data[17686] <= r_data[17685];
                
                r_data[17687] <= r_data[17686];
                
                r_data[17688] <= r_data[17687];
                
                r_data[17689] <= r_data[17688];
                
                r_data[17690] <= r_data[17689];
                
                r_data[17691] <= r_data[17690];
                
                r_data[17692] <= r_data[17691];
                
                r_data[17693] <= r_data[17692];
                
                r_data[17694] <= r_data[17693];
                
                r_data[17695] <= r_data[17694];
                
                r_data[17696] <= r_data[17695];
                
                r_data[17697] <= r_data[17696];
                
                r_data[17698] <= r_data[17697];
                
                r_data[17699] <= r_data[17698];
                
                r_data[17700] <= r_data[17699];
                
                r_data[17701] <= r_data[17700];
                
                r_data[17702] <= r_data[17701];
                
                r_data[17703] <= r_data[17702];
                
                r_data[17704] <= r_data[17703];
                
                r_data[17705] <= r_data[17704];
                
                r_data[17706] <= r_data[17705];
                
                r_data[17707] <= r_data[17706];
                
                r_data[17708] <= r_data[17707];
                
                r_data[17709] <= r_data[17708];
                
                r_data[17710] <= r_data[17709];
                
                r_data[17711] <= r_data[17710];
                
                r_data[17712] <= r_data[17711];
                
                r_data[17713] <= r_data[17712];
                
                r_data[17714] <= r_data[17713];
                
                r_data[17715] <= r_data[17714];
                
                r_data[17716] <= r_data[17715];
                
                r_data[17717] <= r_data[17716];
                
                r_data[17718] <= r_data[17717];
                
                r_data[17719] <= r_data[17718];
                
                r_data[17720] <= r_data[17719];
                
                r_data[17721] <= r_data[17720];
                
                r_data[17722] <= r_data[17721];
                
                r_data[17723] <= r_data[17722];
                
                r_data[17724] <= r_data[17723];
                
                r_data[17725] <= r_data[17724];
                
                r_data[17726] <= r_data[17725];
                
                r_data[17727] <= r_data[17726];
                
                r_data[17728] <= r_data[17727];
                
                r_data[17729] <= r_data[17728];
                
                r_data[17730] <= r_data[17729];
                
                r_data[17731] <= r_data[17730];
                
                r_data[17732] <= r_data[17731];
                
                r_data[17733] <= r_data[17732];
                
                r_data[17734] <= r_data[17733];
                
                r_data[17735] <= r_data[17734];
                
                r_data[17736] <= r_data[17735];
                
                r_data[17737] <= r_data[17736];
                
                r_data[17738] <= r_data[17737];
                
                r_data[17739] <= r_data[17738];
                
                r_data[17740] <= r_data[17739];
                
                r_data[17741] <= r_data[17740];
                
                r_data[17742] <= r_data[17741];
                
                r_data[17743] <= r_data[17742];
                
                r_data[17744] <= r_data[17743];
                
                r_data[17745] <= r_data[17744];
                
                r_data[17746] <= r_data[17745];
                
                r_data[17747] <= r_data[17746];
                
                r_data[17748] <= r_data[17747];
                
                r_data[17749] <= r_data[17748];
                
                r_data[17750] <= r_data[17749];
                
                r_data[17751] <= r_data[17750];
                
                r_data[17752] <= r_data[17751];
                
                r_data[17753] <= r_data[17752];
                
                r_data[17754] <= r_data[17753];
                
                r_data[17755] <= r_data[17754];
                
                r_data[17756] <= r_data[17755];
                
                r_data[17757] <= r_data[17756];
                
                r_data[17758] <= r_data[17757];
                
                r_data[17759] <= r_data[17758];
                
                r_data[17760] <= r_data[17759];
                
                r_data[17761] <= r_data[17760];
                
                r_data[17762] <= r_data[17761];
                
                r_data[17763] <= r_data[17762];
                
                r_data[17764] <= r_data[17763];
                
                r_data[17765] <= r_data[17764];
                
                r_data[17766] <= r_data[17765];
                
                r_data[17767] <= r_data[17766];
                
                r_data[17768] <= r_data[17767];
                
                r_data[17769] <= r_data[17768];
                
                r_data[17770] <= r_data[17769];
                
                r_data[17771] <= r_data[17770];
                
                r_data[17772] <= r_data[17771];
                
                r_data[17773] <= r_data[17772];
                
                r_data[17774] <= r_data[17773];
                
                r_data[17775] <= r_data[17774];
                
                r_data[17776] <= r_data[17775];
                
                r_data[17777] <= r_data[17776];
                
                r_data[17778] <= r_data[17777];
                
                r_data[17779] <= r_data[17778];
                
                r_data[17780] <= r_data[17779];
                
                r_data[17781] <= r_data[17780];
                
                r_data[17782] <= r_data[17781];
                
                r_data[17783] <= r_data[17782];
                
                r_data[17784] <= r_data[17783];
                
                r_data[17785] <= r_data[17784];
                
                r_data[17786] <= r_data[17785];
                
                r_data[17787] <= r_data[17786];
                
                r_data[17788] <= r_data[17787];
                
                r_data[17789] <= r_data[17788];
                
                r_data[17790] <= r_data[17789];
                
                r_data[17791] <= r_data[17790];
                
                r_data[17792] <= r_data[17791];
                
                r_data[17793] <= r_data[17792];
                
                r_data[17794] <= r_data[17793];
                
                r_data[17795] <= r_data[17794];
                
                r_data[17796] <= r_data[17795];
                
                r_data[17797] <= r_data[17796];
                
                r_data[17798] <= r_data[17797];
                
                r_data[17799] <= r_data[17798];
                
                r_data[17800] <= r_data[17799];
                
                r_data[17801] <= r_data[17800];
                
                r_data[17802] <= r_data[17801];
                
                r_data[17803] <= r_data[17802];
                
                r_data[17804] <= r_data[17803];
                
                r_data[17805] <= r_data[17804];
                
                r_data[17806] <= r_data[17805];
                
                r_data[17807] <= r_data[17806];
                
                r_data[17808] <= r_data[17807];
                
                r_data[17809] <= r_data[17808];
                
                r_data[17810] <= r_data[17809];
                
                r_data[17811] <= r_data[17810];
                
                r_data[17812] <= r_data[17811];
                
                r_data[17813] <= r_data[17812];
                
                r_data[17814] <= r_data[17813];
                
                r_data[17815] <= r_data[17814];
                
                r_data[17816] <= r_data[17815];
                
                r_data[17817] <= r_data[17816];
                
                r_data[17818] <= r_data[17817];
                
                r_data[17819] <= r_data[17818];
                
                r_data[17820] <= r_data[17819];
                
                r_data[17821] <= r_data[17820];
                
                r_data[17822] <= r_data[17821];
                
                r_data[17823] <= r_data[17822];
                
                r_data[17824] <= r_data[17823];
                
                r_data[17825] <= r_data[17824];
                
                r_data[17826] <= r_data[17825];
                
                r_data[17827] <= r_data[17826];
                
                r_data[17828] <= r_data[17827];
                
                r_data[17829] <= r_data[17828];
                
                r_data[17830] <= r_data[17829];
                
                r_data[17831] <= r_data[17830];
                
                r_data[17832] <= r_data[17831];
                
                r_data[17833] <= r_data[17832];
                
                r_data[17834] <= r_data[17833];
                
                r_data[17835] <= r_data[17834];
                
                r_data[17836] <= r_data[17835];
                
                r_data[17837] <= r_data[17836];
                
                r_data[17838] <= r_data[17837];
                
                r_data[17839] <= r_data[17838];
                
                r_data[17840] <= r_data[17839];
                
                r_data[17841] <= r_data[17840];
                
                r_data[17842] <= r_data[17841];
                
                r_data[17843] <= r_data[17842];
                
                r_data[17844] <= r_data[17843];
                
                r_data[17845] <= r_data[17844];
                
                r_data[17846] <= r_data[17845];
                
                r_data[17847] <= r_data[17846];
                
                r_data[17848] <= r_data[17847];
                
                r_data[17849] <= r_data[17848];
                
                r_data[17850] <= r_data[17849];
                
                r_data[17851] <= r_data[17850];
                
                r_data[17852] <= r_data[17851];
                
                r_data[17853] <= r_data[17852];
                
                r_data[17854] <= r_data[17853];
                
                r_data[17855] <= r_data[17854];
                
                r_data[17856] <= r_data[17855];
                
                r_data[17857] <= r_data[17856];
                
                r_data[17858] <= r_data[17857];
                
                r_data[17859] <= r_data[17858];
                
                r_data[17860] <= r_data[17859];
                
                r_data[17861] <= r_data[17860];
                
                r_data[17862] <= r_data[17861];
                
                r_data[17863] <= r_data[17862];
                
                r_data[17864] <= r_data[17863];
                
                r_data[17865] <= r_data[17864];
                
                r_data[17866] <= r_data[17865];
                
                r_data[17867] <= r_data[17866];
                
                r_data[17868] <= r_data[17867];
                
                r_data[17869] <= r_data[17868];
                
                r_data[17870] <= r_data[17869];
                
                r_data[17871] <= r_data[17870];
                
                r_data[17872] <= r_data[17871];
                
                r_data[17873] <= r_data[17872];
                
                r_data[17874] <= r_data[17873];
                
                r_data[17875] <= r_data[17874];
                
                r_data[17876] <= r_data[17875];
                
                r_data[17877] <= r_data[17876];
                
                r_data[17878] <= r_data[17877];
                
                r_data[17879] <= r_data[17878];
                
                r_data[17880] <= r_data[17879];
                
                r_data[17881] <= r_data[17880];
                
                r_data[17882] <= r_data[17881];
                
                r_data[17883] <= r_data[17882];
                
                r_data[17884] <= r_data[17883];
                
                r_data[17885] <= r_data[17884];
                
                r_data[17886] <= r_data[17885];
                
                r_data[17887] <= r_data[17886];
                
                r_data[17888] <= r_data[17887];
                
                r_data[17889] <= r_data[17888];
                
                r_data[17890] <= r_data[17889];
                
                r_data[17891] <= r_data[17890];
                
                r_data[17892] <= r_data[17891];
                
                r_data[17893] <= r_data[17892];
                
                r_data[17894] <= r_data[17893];
                
                r_data[17895] <= r_data[17894];
                
                r_data[17896] <= r_data[17895];
                
                r_data[17897] <= r_data[17896];
                
                r_data[17898] <= r_data[17897];
                
                r_data[17899] <= r_data[17898];
                
                r_data[17900] <= r_data[17899];
                
                r_data[17901] <= r_data[17900];
                
                r_data[17902] <= r_data[17901];
                
                r_data[17903] <= r_data[17902];
                
                r_data[17904] <= r_data[17903];
                
                r_data[17905] <= r_data[17904];
                
                r_data[17906] <= r_data[17905];
                
                r_data[17907] <= r_data[17906];
                
                r_data[17908] <= r_data[17907];
                
                r_data[17909] <= r_data[17908];
                
                r_data[17910] <= r_data[17909];
                
                r_data[17911] <= r_data[17910];
                
                r_data[17912] <= r_data[17911];
                
                r_data[17913] <= r_data[17912];
                
                r_data[17914] <= r_data[17913];
                
                r_data[17915] <= r_data[17914];
                
                r_data[17916] <= r_data[17915];
                
                r_data[17917] <= r_data[17916];
                
                r_data[17918] <= r_data[17917];
                
                r_data[17919] <= r_data[17918];
                
                r_data[17920] <= r_data[17919];
                
                r_data[17921] <= r_data[17920];
                
                r_data[17922] <= r_data[17921];
                
                r_data[17923] <= r_data[17922];
                
                r_data[17924] <= r_data[17923];
                
                r_data[17925] <= r_data[17924];
                
                r_data[17926] <= r_data[17925];
                
                r_data[17927] <= r_data[17926];
                
                r_data[17928] <= r_data[17927];
                
                r_data[17929] <= r_data[17928];
                
                r_data[17930] <= r_data[17929];
                
                r_data[17931] <= r_data[17930];
                
                r_data[17932] <= r_data[17931];
                
                r_data[17933] <= r_data[17932];
                
                r_data[17934] <= r_data[17933];
                
                r_data[17935] <= r_data[17934];
                
                r_data[17936] <= r_data[17935];
                
                r_data[17937] <= r_data[17936];
                
                r_data[17938] <= r_data[17937];
                
                r_data[17939] <= r_data[17938];
                
                r_data[17940] <= r_data[17939];
                
                r_data[17941] <= r_data[17940];
                
                r_data[17942] <= r_data[17941];
                
                r_data[17943] <= r_data[17942];
                
                r_data[17944] <= r_data[17943];
                
                r_data[17945] <= r_data[17944];
                
                r_data[17946] <= r_data[17945];
                
                r_data[17947] <= r_data[17946];
                
                r_data[17948] <= r_data[17947];
                
                r_data[17949] <= r_data[17948];
                
                r_data[17950] <= r_data[17949];
                
                r_data[17951] <= r_data[17950];
                
                r_data[17952] <= r_data[17951];
                
                r_data[17953] <= r_data[17952];
                
                r_data[17954] <= r_data[17953];
                
                r_data[17955] <= r_data[17954];
                
                r_data[17956] <= r_data[17955];
                
                r_data[17957] <= r_data[17956];
                
                r_data[17958] <= r_data[17957];
                
                r_data[17959] <= r_data[17958];
                
                r_data[17960] <= r_data[17959];
                
                r_data[17961] <= r_data[17960];
                
                r_data[17962] <= r_data[17961];
                
                r_data[17963] <= r_data[17962];
                
                r_data[17964] <= r_data[17963];
                
                r_data[17965] <= r_data[17964];
                
                r_data[17966] <= r_data[17965];
                
                r_data[17967] <= r_data[17966];
                
                r_data[17968] <= r_data[17967];
                
                r_data[17969] <= r_data[17968];
                
                r_data[17970] <= r_data[17969];
                
                r_data[17971] <= r_data[17970];
                
                r_data[17972] <= r_data[17971];
                
                r_data[17973] <= r_data[17972];
                
                r_data[17974] <= r_data[17973];
                
                r_data[17975] <= r_data[17974];
                
                r_data[17976] <= r_data[17975];
                
                r_data[17977] <= r_data[17976];
                
                r_data[17978] <= r_data[17977];
                
                r_data[17979] <= r_data[17978];
                
                r_data[17980] <= r_data[17979];
                
                r_data[17981] <= r_data[17980];
                
                r_data[17982] <= r_data[17981];
                
                r_data[17983] <= r_data[17982];
                
                r_data[17984] <= r_data[17983];
                
                r_data[17985] <= r_data[17984];
                
                r_data[17986] <= r_data[17985];
                
                r_data[17987] <= r_data[17986];
                
                r_data[17988] <= r_data[17987];
                
                r_data[17989] <= r_data[17988];
                
                r_data[17990] <= r_data[17989];
                
                r_data[17991] <= r_data[17990];
                
                r_data[17992] <= r_data[17991];
                
                r_data[17993] <= r_data[17992];
                
                r_data[17994] <= r_data[17993];
                
                r_data[17995] <= r_data[17994];
                
                r_data[17996] <= r_data[17995];
                
                r_data[17997] <= r_data[17996];
                
                r_data[17998] <= r_data[17997];
                
                r_data[17999] <= r_data[17998];
                
                r_data[18000] <= r_data[17999];
                
                r_data[18001] <= r_data[18000];
                
                r_data[18002] <= r_data[18001];
                
                r_data[18003] <= r_data[18002];
                
                r_data[18004] <= r_data[18003];
                
                r_data[18005] <= r_data[18004];
                
                r_data[18006] <= r_data[18005];
                
                r_data[18007] <= r_data[18006];
                
                r_data[18008] <= r_data[18007];
                
                r_data[18009] <= r_data[18008];
                
                r_data[18010] <= r_data[18009];
                
                r_data[18011] <= r_data[18010];
                
                r_data[18012] <= r_data[18011];
                
                r_data[18013] <= r_data[18012];
                
                r_data[18014] <= r_data[18013];
                
                r_data[18015] <= r_data[18014];
                
                r_data[18016] <= r_data[18015];
                
                r_data[18017] <= r_data[18016];
                
                r_data[18018] <= r_data[18017];
                
                r_data[18019] <= r_data[18018];
                
                r_data[18020] <= r_data[18019];
                
                r_data[18021] <= r_data[18020];
                
                r_data[18022] <= r_data[18021];
                
                r_data[18023] <= r_data[18022];
                
                r_data[18024] <= r_data[18023];
                
                r_data[18025] <= r_data[18024];
                
                r_data[18026] <= r_data[18025];
                
                r_data[18027] <= r_data[18026];
                
                r_data[18028] <= r_data[18027];
                
                r_data[18029] <= r_data[18028];
                
                r_data[18030] <= r_data[18029];
                
                r_data[18031] <= r_data[18030];
                
                r_data[18032] <= r_data[18031];
                
                r_data[18033] <= r_data[18032];
                
                r_data[18034] <= r_data[18033];
                
                r_data[18035] <= r_data[18034];
                
                r_data[18036] <= r_data[18035];
                
                r_data[18037] <= r_data[18036];
                
                r_data[18038] <= r_data[18037];
                
                r_data[18039] <= r_data[18038];
                
                r_data[18040] <= r_data[18039];
                
                r_data[18041] <= r_data[18040];
                
                r_data[18042] <= r_data[18041];
                
                r_data[18043] <= r_data[18042];
                
                r_data[18044] <= r_data[18043];
                
                r_data[18045] <= r_data[18044];
                
                r_data[18046] <= r_data[18045];
                
                r_data[18047] <= r_data[18046];
                
                r_data[18048] <= r_data[18047];
                
                r_data[18049] <= r_data[18048];
                
                r_data[18050] <= r_data[18049];
                
                r_data[18051] <= r_data[18050];
                
                r_data[18052] <= r_data[18051];
                
                r_data[18053] <= r_data[18052];
                
                r_data[18054] <= r_data[18053];
                
                r_data[18055] <= r_data[18054];
                
                r_data[18056] <= r_data[18055];
                
                r_data[18057] <= r_data[18056];
                
                r_data[18058] <= r_data[18057];
                
                r_data[18059] <= r_data[18058];
                
                r_data[18060] <= r_data[18059];
                
                r_data[18061] <= r_data[18060];
                
                r_data[18062] <= r_data[18061];
                
                r_data[18063] <= r_data[18062];
                
                r_data[18064] <= r_data[18063];
                
                r_data[18065] <= r_data[18064];
                
                r_data[18066] <= r_data[18065];
                
                r_data[18067] <= r_data[18066];
                
                r_data[18068] <= r_data[18067];
                
                r_data[18069] <= r_data[18068];
                
                r_data[18070] <= r_data[18069];
                
                r_data[18071] <= r_data[18070];
                
                r_data[18072] <= r_data[18071];
                
                r_data[18073] <= r_data[18072];
                
                r_data[18074] <= r_data[18073];
                
                r_data[18075] <= r_data[18074];
                
                r_data[18076] <= r_data[18075];
                
                r_data[18077] <= r_data[18076];
                
                r_data[18078] <= r_data[18077];
                
                r_data[18079] <= r_data[18078];
                
                r_data[18080] <= r_data[18079];
                
                r_data[18081] <= r_data[18080];
                
                r_data[18082] <= r_data[18081];
                
                r_data[18083] <= r_data[18082];
                
                r_data[18084] <= r_data[18083];
                
                r_data[18085] <= r_data[18084];
                
                r_data[18086] <= r_data[18085];
                
                r_data[18087] <= r_data[18086];
                
                r_data[18088] <= r_data[18087];
                
                r_data[18089] <= r_data[18088];
                
                r_data[18090] <= r_data[18089];
                
                r_data[18091] <= r_data[18090];
                
                r_data[18092] <= r_data[18091];
                
                r_data[18093] <= r_data[18092];
                
                r_data[18094] <= r_data[18093];
                
                r_data[18095] <= r_data[18094];
                
                r_data[18096] <= r_data[18095];
                
                r_data[18097] <= r_data[18096];
                
                r_data[18098] <= r_data[18097];
                
                r_data[18099] <= r_data[18098];
                
                r_data[18100] <= r_data[18099];
                
                r_data[18101] <= r_data[18100];
                
                r_data[18102] <= r_data[18101];
                
                r_data[18103] <= r_data[18102];
                
                r_data[18104] <= r_data[18103];
                
                r_data[18105] <= r_data[18104];
                
                r_data[18106] <= r_data[18105];
                
                r_data[18107] <= r_data[18106];
                
                r_data[18108] <= r_data[18107];
                
                r_data[18109] <= r_data[18108];
                
                r_data[18110] <= r_data[18109];
                
                r_data[18111] <= r_data[18110];
                
                r_data[18112] <= r_data[18111];
                
                r_data[18113] <= r_data[18112];
                
                r_data[18114] <= r_data[18113];
                
                r_data[18115] <= r_data[18114];
                
                r_data[18116] <= r_data[18115];
                
                r_data[18117] <= r_data[18116];
                
                r_data[18118] <= r_data[18117];
                
                r_data[18119] <= r_data[18118];
                
                r_data[18120] <= r_data[18119];
                
                r_data[18121] <= r_data[18120];
                
                r_data[18122] <= r_data[18121];
                
                r_data[18123] <= r_data[18122];
                
                r_data[18124] <= r_data[18123];
                
                r_data[18125] <= r_data[18124];
                
                r_data[18126] <= r_data[18125];
                
                r_data[18127] <= r_data[18126];
                
                r_data[18128] <= r_data[18127];
                
                r_data[18129] <= r_data[18128];
                
                r_data[18130] <= r_data[18129];
                
                r_data[18131] <= r_data[18130];
                
                r_data[18132] <= r_data[18131];
                
                r_data[18133] <= r_data[18132];
                
                r_data[18134] <= r_data[18133];
                
                r_data[18135] <= r_data[18134];
                
                r_data[18136] <= r_data[18135];
                
                r_data[18137] <= r_data[18136];
                
                r_data[18138] <= r_data[18137];
                
                r_data[18139] <= r_data[18138];
                
                r_data[18140] <= r_data[18139];
                
                r_data[18141] <= r_data[18140];
                
                r_data[18142] <= r_data[18141];
                
                r_data[18143] <= r_data[18142];
                
                r_data[18144] <= r_data[18143];
                
                r_data[18145] <= r_data[18144];
                
                r_data[18146] <= r_data[18145];
                
                r_data[18147] <= r_data[18146];
                
                r_data[18148] <= r_data[18147];
                
                r_data[18149] <= r_data[18148];
                
                r_data[18150] <= r_data[18149];
                
                r_data[18151] <= r_data[18150];
                
                r_data[18152] <= r_data[18151];
                
                r_data[18153] <= r_data[18152];
                
                r_data[18154] <= r_data[18153];
                
                r_data[18155] <= r_data[18154];
                
                r_data[18156] <= r_data[18155];
                
                r_data[18157] <= r_data[18156];
                
                r_data[18158] <= r_data[18157];
                
                r_data[18159] <= r_data[18158];
                
                r_data[18160] <= r_data[18159];
                
                r_data[18161] <= r_data[18160];
                
                r_data[18162] <= r_data[18161];
                
                r_data[18163] <= r_data[18162];
                
                r_data[18164] <= r_data[18163];
                
                r_data[18165] <= r_data[18164];
                
                r_data[18166] <= r_data[18165];
                
                r_data[18167] <= r_data[18166];
                
                r_data[18168] <= r_data[18167];
                
                r_data[18169] <= r_data[18168];
                
                r_data[18170] <= r_data[18169];
                
                r_data[18171] <= r_data[18170];
                
                r_data[18172] <= r_data[18171];
                
                r_data[18173] <= r_data[18172];
                
                r_data[18174] <= r_data[18173];
                
                r_data[18175] <= r_data[18174];
                
                r_data[18176] <= r_data[18175];
                
                r_data[18177] <= r_data[18176];
                
                r_data[18178] <= r_data[18177];
                
                r_data[18179] <= r_data[18178];
                
                r_data[18180] <= r_data[18179];
                
                r_data[18181] <= r_data[18180];
                
                r_data[18182] <= r_data[18181];
                
                r_data[18183] <= r_data[18182];
                
                r_data[18184] <= r_data[18183];
                
                r_data[18185] <= r_data[18184];
                
                r_data[18186] <= r_data[18185];
                
                r_data[18187] <= r_data[18186];
                
                r_data[18188] <= r_data[18187];
                
                r_data[18189] <= r_data[18188];
                
                r_data[18190] <= r_data[18189];
                
                r_data[18191] <= r_data[18190];
                
                r_data[18192] <= r_data[18191];
                
                r_data[18193] <= r_data[18192];
                
                r_data[18194] <= r_data[18193];
                
                r_data[18195] <= r_data[18194];
                
                r_data[18196] <= r_data[18195];
                
                r_data[18197] <= r_data[18196];
                
                r_data[18198] <= r_data[18197];
                
                r_data[18199] <= r_data[18198];
                
                r_data[18200] <= r_data[18199];
                
                r_data[18201] <= r_data[18200];
                
                r_data[18202] <= r_data[18201];
                
                r_data[18203] <= r_data[18202];
                
                r_data[18204] <= r_data[18203];
                
                r_data[18205] <= r_data[18204];
                
                r_data[18206] <= r_data[18205];
                
                r_data[18207] <= r_data[18206];
                
                r_data[18208] <= r_data[18207];
                
                r_data[18209] <= r_data[18208];
                
                r_data[18210] <= r_data[18209];
                
                r_data[18211] <= r_data[18210];
                
                r_data[18212] <= r_data[18211];
                
                r_data[18213] <= r_data[18212];
                
                r_data[18214] <= r_data[18213];
                
                r_data[18215] <= r_data[18214];
                
                r_data[18216] <= r_data[18215];
                
                r_data[18217] <= r_data[18216];
                
                r_data[18218] <= r_data[18217];
                
                r_data[18219] <= r_data[18218];
                
                r_data[18220] <= r_data[18219];
                
                r_data[18221] <= r_data[18220];
                
                r_data[18222] <= r_data[18221];
                
                r_data[18223] <= r_data[18222];
                
                r_data[18224] <= r_data[18223];
                
                r_data[18225] <= r_data[18224];
                
                r_data[18226] <= r_data[18225];
                
                r_data[18227] <= r_data[18226];
                
                r_data[18228] <= r_data[18227];
                
                r_data[18229] <= r_data[18228];
                
                r_data[18230] <= r_data[18229];
                
                r_data[18231] <= r_data[18230];
                
                r_data[18232] <= r_data[18231];
                
                r_data[18233] <= r_data[18232];
                
                r_data[18234] <= r_data[18233];
                
                r_data[18235] <= r_data[18234];
                
                r_data[18236] <= r_data[18235];
                
                r_data[18237] <= r_data[18236];
                
                r_data[18238] <= r_data[18237];
                
                r_data[18239] <= r_data[18238];
                
                r_data[18240] <= r_data[18239];
                
                r_data[18241] <= r_data[18240];
                
                r_data[18242] <= r_data[18241];
                
                r_data[18243] <= r_data[18242];
                
                r_data[18244] <= r_data[18243];
                
                r_data[18245] <= r_data[18244];
                
                r_data[18246] <= r_data[18245];
                
                r_data[18247] <= r_data[18246];
                
                r_data[18248] <= r_data[18247];
                
                r_data[18249] <= r_data[18248];
                
                r_data[18250] <= r_data[18249];
                
                r_data[18251] <= r_data[18250];
                
                r_data[18252] <= r_data[18251];
                
                r_data[18253] <= r_data[18252];
                
                r_data[18254] <= r_data[18253];
                
                r_data[18255] <= r_data[18254];
                
                r_data[18256] <= r_data[18255];
                
                r_data[18257] <= r_data[18256];
                
                r_data[18258] <= r_data[18257];
                
                r_data[18259] <= r_data[18258];
                
                r_data[18260] <= r_data[18259];
                
                r_data[18261] <= r_data[18260];
                
                r_data[18262] <= r_data[18261];
                
                r_data[18263] <= r_data[18262];
                
                r_data[18264] <= r_data[18263];
                
                r_data[18265] <= r_data[18264];
                
                r_data[18266] <= r_data[18265];
                
                r_data[18267] <= r_data[18266];
                
                r_data[18268] <= r_data[18267];
                
                r_data[18269] <= r_data[18268];
                
                r_data[18270] <= r_data[18269];
                
                r_data[18271] <= r_data[18270];
                
                r_data[18272] <= r_data[18271];
                
                r_data[18273] <= r_data[18272];
                
                r_data[18274] <= r_data[18273];
                
                r_data[18275] <= r_data[18274];
                
                r_data[18276] <= r_data[18275];
                
                r_data[18277] <= r_data[18276];
                
                r_data[18278] <= r_data[18277];
                
                r_data[18279] <= r_data[18278];
                
                r_data[18280] <= r_data[18279];
                
                r_data[18281] <= r_data[18280];
                
                r_data[18282] <= r_data[18281];
                
                r_data[18283] <= r_data[18282];
                
                r_data[18284] <= r_data[18283];
                
                r_data[18285] <= r_data[18284];
                
                r_data[18286] <= r_data[18285];
                
                r_data[18287] <= r_data[18286];
                
                r_data[18288] <= r_data[18287];
                
                r_data[18289] <= r_data[18288];
                
                r_data[18290] <= r_data[18289];
                
                r_data[18291] <= r_data[18290];
                
                r_data[18292] <= r_data[18291];
                
                r_data[18293] <= r_data[18292];
                
                r_data[18294] <= r_data[18293];
                
                r_data[18295] <= r_data[18294];
                
                r_data[18296] <= r_data[18295];
                
                r_data[18297] <= r_data[18296];
                
                r_data[18298] <= r_data[18297];
                
                r_data[18299] <= r_data[18298];
                
                r_data[18300] <= r_data[18299];
                
                r_data[18301] <= r_data[18300];
                
                r_data[18302] <= r_data[18301];
                
                r_data[18303] <= r_data[18302];
                
                r_data[18304] <= r_data[18303];
                
                r_data[18305] <= r_data[18304];
                
                r_data[18306] <= r_data[18305];
                
                r_data[18307] <= r_data[18306];
                
                r_data[18308] <= r_data[18307];
                
                r_data[18309] <= r_data[18308];
                
                r_data[18310] <= r_data[18309];
                
                r_data[18311] <= r_data[18310];
                
                r_data[18312] <= r_data[18311];
                
                r_data[18313] <= r_data[18312];
                
                r_data[18314] <= r_data[18313];
                
                r_data[18315] <= r_data[18314];
                
                r_data[18316] <= r_data[18315];
                
                r_data[18317] <= r_data[18316];
                
                r_data[18318] <= r_data[18317];
                
                r_data[18319] <= r_data[18318];
                
                r_data[18320] <= r_data[18319];
                
                r_data[18321] <= r_data[18320];
                
                r_data[18322] <= r_data[18321];
                
                r_data[18323] <= r_data[18322];
                
                r_data[18324] <= r_data[18323];
                
                r_data[18325] <= r_data[18324];
                
                r_data[18326] <= r_data[18325];
                
                r_data[18327] <= r_data[18326];
                
                r_data[18328] <= r_data[18327];
                
                r_data[18329] <= r_data[18328];
                
                r_data[18330] <= r_data[18329];
                
                r_data[18331] <= r_data[18330];
                
                r_data[18332] <= r_data[18331];
                
                r_data[18333] <= r_data[18332];
                
                r_data[18334] <= r_data[18333];
                
                r_data[18335] <= r_data[18334];
                
                r_data[18336] <= r_data[18335];
                
                r_data[18337] <= r_data[18336];
                
                r_data[18338] <= r_data[18337];
                
                r_data[18339] <= r_data[18338];
                
                r_data[18340] <= r_data[18339];
                
                r_data[18341] <= r_data[18340];
                
                r_data[18342] <= r_data[18341];
                
                r_data[18343] <= r_data[18342];
                
                r_data[18344] <= r_data[18343];
                
                r_data[18345] <= r_data[18344];
                
                r_data[18346] <= r_data[18345];
                
                r_data[18347] <= r_data[18346];
                
                r_data[18348] <= r_data[18347];
                
                r_data[18349] <= r_data[18348];
                
                r_data[18350] <= r_data[18349];
                
                r_data[18351] <= r_data[18350];
                
                r_data[18352] <= r_data[18351];
                
                r_data[18353] <= r_data[18352];
                
                r_data[18354] <= r_data[18353];
                
                r_data[18355] <= r_data[18354];
                
                r_data[18356] <= r_data[18355];
                
                r_data[18357] <= r_data[18356];
                
                r_data[18358] <= r_data[18357];
                
                r_data[18359] <= r_data[18358];
                
                r_data[18360] <= r_data[18359];
                
                r_data[18361] <= r_data[18360];
                
                r_data[18362] <= r_data[18361];
                
                r_data[18363] <= r_data[18362];
                
                r_data[18364] <= r_data[18363];
                
                r_data[18365] <= r_data[18364];
                
                r_data[18366] <= r_data[18365];
                
                r_data[18367] <= r_data[18366];
                
                r_data[18368] <= r_data[18367];
                
                r_data[18369] <= r_data[18368];
                
                r_data[18370] <= r_data[18369];
                
                r_data[18371] <= r_data[18370];
                
                r_data[18372] <= r_data[18371];
                
                r_data[18373] <= r_data[18372];
                
                r_data[18374] <= r_data[18373];
                
                r_data[18375] <= r_data[18374];
                
                r_data[18376] <= r_data[18375];
                
                r_data[18377] <= r_data[18376];
                
                r_data[18378] <= r_data[18377];
                
                r_data[18379] <= r_data[18378];
                
                r_data[18380] <= r_data[18379];
                
                r_data[18381] <= r_data[18380];
                
                r_data[18382] <= r_data[18381];
                
                r_data[18383] <= r_data[18382];
                
                r_data[18384] <= r_data[18383];
                
                r_data[18385] <= r_data[18384];
                
                r_data[18386] <= r_data[18385];
                
                r_data[18387] <= r_data[18386];
                
                r_data[18388] <= r_data[18387];
                
                r_data[18389] <= r_data[18388];
                
                r_data[18390] <= r_data[18389];
                
                r_data[18391] <= r_data[18390];
                
                r_data[18392] <= r_data[18391];
                
                r_data[18393] <= r_data[18392];
                
                r_data[18394] <= r_data[18393];
                
                r_data[18395] <= r_data[18394];
                
                r_data[18396] <= r_data[18395];
                
                r_data[18397] <= r_data[18396];
                
                r_data[18398] <= r_data[18397];
                
                r_data[18399] <= r_data[18398];
                
                r_data[18400] <= r_data[18399];
                
                r_data[18401] <= r_data[18400];
                
                r_data[18402] <= r_data[18401];
                
                r_data[18403] <= r_data[18402];
                
                r_data[18404] <= r_data[18403];
                
                r_data[18405] <= r_data[18404];
                
                r_data[18406] <= r_data[18405];
                
                r_data[18407] <= r_data[18406];
                
                r_data[18408] <= r_data[18407];
                
                r_data[18409] <= r_data[18408];
                
                r_data[18410] <= r_data[18409];
                
                r_data[18411] <= r_data[18410];
                
                r_data[18412] <= r_data[18411];
                
                r_data[18413] <= r_data[18412];
                
                r_data[18414] <= r_data[18413];
                
                r_data[18415] <= r_data[18414];
                
                r_data[18416] <= r_data[18415];
                
                r_data[18417] <= r_data[18416];
                
                r_data[18418] <= r_data[18417];
                
                r_data[18419] <= r_data[18418];
                
                r_data[18420] <= r_data[18419];
                
                r_data[18421] <= r_data[18420];
                
                r_data[18422] <= r_data[18421];
                
                r_data[18423] <= r_data[18422];
                
                r_data[18424] <= r_data[18423];
                
                r_data[18425] <= r_data[18424];
                
                r_data[18426] <= r_data[18425];
                
                r_data[18427] <= r_data[18426];
                
                r_data[18428] <= r_data[18427];
                
                r_data[18429] <= r_data[18428];
                
                r_data[18430] <= r_data[18429];
                
                r_data[18431] <= r_data[18430];
                
                r_data[18432] <= r_data[18431];
                
                r_data[18433] <= r_data[18432];
                
                r_data[18434] <= r_data[18433];
                
                r_data[18435] <= r_data[18434];
                
                r_data[18436] <= r_data[18435];
                
                r_data[18437] <= r_data[18436];
                
                r_data[18438] <= r_data[18437];
                
                r_data[18439] <= r_data[18438];
                
                r_data[18440] <= r_data[18439];
                
                r_data[18441] <= r_data[18440];
                
                r_data[18442] <= r_data[18441];
                
                r_data[18443] <= r_data[18442];
                
                r_data[18444] <= r_data[18443];
                
                r_data[18445] <= r_data[18444];
                
                r_data[18446] <= r_data[18445];
                
                r_data[18447] <= r_data[18446];
                
                r_data[18448] <= r_data[18447];
                
                r_data[18449] <= r_data[18448];
                
                r_data[18450] <= r_data[18449];
                
                r_data[18451] <= r_data[18450];
                
                r_data[18452] <= r_data[18451];
                
                r_data[18453] <= r_data[18452];
                
                r_data[18454] <= r_data[18453];
                
                r_data[18455] <= r_data[18454];
                
                r_data[18456] <= r_data[18455];
                
                r_data[18457] <= r_data[18456];
                
                r_data[18458] <= r_data[18457];
                
                r_data[18459] <= r_data[18458];
                
                r_data[18460] <= r_data[18459];
                
                r_data[18461] <= r_data[18460];
                
                r_data[18462] <= r_data[18461];
                
                r_data[18463] <= r_data[18462];
                
                r_data[18464] <= r_data[18463];
                
                r_data[18465] <= r_data[18464];
                
                r_data[18466] <= r_data[18465];
                
                r_data[18467] <= r_data[18466];
                
                r_data[18468] <= r_data[18467];
                
                r_data[18469] <= r_data[18468];
                
                r_data[18470] <= r_data[18469];
                
                r_data[18471] <= r_data[18470];
                
                r_data[18472] <= r_data[18471];
                
                r_data[18473] <= r_data[18472];
                
                r_data[18474] <= r_data[18473];
                
                r_data[18475] <= r_data[18474];
                
                r_data[18476] <= r_data[18475];
                
                r_data[18477] <= r_data[18476];
                
                r_data[18478] <= r_data[18477];
                
                r_data[18479] <= r_data[18478];
                
                r_data[18480] <= r_data[18479];
                
                r_data[18481] <= r_data[18480];
                
                r_data[18482] <= r_data[18481];
                
                r_data[18483] <= r_data[18482];
                
                r_data[18484] <= r_data[18483];
                
                r_data[18485] <= r_data[18484];
                
                r_data[18486] <= r_data[18485];
                
                r_data[18487] <= r_data[18486];
                
                r_data[18488] <= r_data[18487];
                
                r_data[18489] <= r_data[18488];
                
                r_data[18490] <= r_data[18489];
                
                r_data[18491] <= r_data[18490];
                
                r_data[18492] <= r_data[18491];
                
                r_data[18493] <= r_data[18492];
                
                r_data[18494] <= r_data[18493];
                
                r_data[18495] <= r_data[18494];
                
                r_data[18496] <= r_data[18495];
                
                r_data[18497] <= r_data[18496];
                
                r_data[18498] <= r_data[18497];
                
                r_data[18499] <= r_data[18498];
                
                r_data[18500] <= r_data[18499];
                
                r_data[18501] <= r_data[18500];
                
                r_data[18502] <= r_data[18501];
                
                r_data[18503] <= r_data[18502];
                
                r_data[18504] <= r_data[18503];
                
                r_data[18505] <= r_data[18504];
                
                r_data[18506] <= r_data[18505];
                
                r_data[18507] <= r_data[18506];
                
                r_data[18508] <= r_data[18507];
                
                r_data[18509] <= r_data[18508];
                
                r_data[18510] <= r_data[18509];
                
                r_data[18511] <= r_data[18510];
                
                r_data[18512] <= r_data[18511];
                
                r_data[18513] <= r_data[18512];
                
                r_data[18514] <= r_data[18513];
                
                r_data[18515] <= r_data[18514];
                
                r_data[18516] <= r_data[18515];
                
                r_data[18517] <= r_data[18516];
                
                r_data[18518] <= r_data[18517];
                
                r_data[18519] <= r_data[18518];
                
                r_data[18520] <= r_data[18519];
                
                r_data[18521] <= r_data[18520];
                
                r_data[18522] <= r_data[18521];
                
                r_data[18523] <= r_data[18522];
                
                r_data[18524] <= r_data[18523];
                
                r_data[18525] <= r_data[18524];
                
                r_data[18526] <= r_data[18525];
                
                r_data[18527] <= r_data[18526];
                
                r_data[18528] <= r_data[18527];
                
                r_data[18529] <= r_data[18528];
                
                r_data[18530] <= r_data[18529];
                
                r_data[18531] <= r_data[18530];
                
                r_data[18532] <= r_data[18531];
                
                r_data[18533] <= r_data[18532];
                
                r_data[18534] <= r_data[18533];
                
                r_data[18535] <= r_data[18534];
                
                r_data[18536] <= r_data[18535];
                
                r_data[18537] <= r_data[18536];
                
                r_data[18538] <= r_data[18537];
                
                r_data[18539] <= r_data[18538];
                
                r_data[18540] <= r_data[18539];
                
                r_data[18541] <= r_data[18540];
                
                r_data[18542] <= r_data[18541];
                
                r_data[18543] <= r_data[18542];
                
                r_data[18544] <= r_data[18543];
                
                r_data[18545] <= r_data[18544];
                
                r_data[18546] <= r_data[18545];
                
                r_data[18547] <= r_data[18546];
                
                r_data[18548] <= r_data[18547];
                
                r_data[18549] <= r_data[18548];
                
                r_data[18550] <= r_data[18549];
                
                r_data[18551] <= r_data[18550];
                
                r_data[18552] <= r_data[18551];
                
                r_data[18553] <= r_data[18552];
                
                r_data[18554] <= r_data[18553];
                
                r_data[18555] <= r_data[18554];
                
                r_data[18556] <= r_data[18555];
                
                r_data[18557] <= r_data[18556];
                
                r_data[18558] <= r_data[18557];
                
                r_data[18559] <= r_data[18558];
                
                r_data[18560] <= r_data[18559];
                
                r_data[18561] <= r_data[18560];
                
                r_data[18562] <= r_data[18561];
                
                r_data[18563] <= r_data[18562];
                
                r_data[18564] <= r_data[18563];
                
                r_data[18565] <= r_data[18564];
                
                r_data[18566] <= r_data[18565];
                
                r_data[18567] <= r_data[18566];
                
                r_data[18568] <= r_data[18567];
                
                r_data[18569] <= r_data[18568];
                
                r_data[18570] <= r_data[18569];
                
                r_data[18571] <= r_data[18570];
                
                r_data[18572] <= r_data[18571];
                
                r_data[18573] <= r_data[18572];
                
                r_data[18574] <= r_data[18573];
                
                r_data[18575] <= r_data[18574];
                
                r_data[18576] <= r_data[18575];
                
                r_data[18577] <= r_data[18576];
                
                r_data[18578] <= r_data[18577];
                
                r_data[18579] <= r_data[18578];
                
                r_data[18580] <= r_data[18579];
                
                r_data[18581] <= r_data[18580];
                
                r_data[18582] <= r_data[18581];
                
                r_data[18583] <= r_data[18582];
                
                r_data[18584] <= r_data[18583];
                
                r_data[18585] <= r_data[18584];
                
                r_data[18586] <= r_data[18585];
                
                r_data[18587] <= r_data[18586];
                
                r_data[18588] <= r_data[18587];
                
                r_data[18589] <= r_data[18588];
                
                r_data[18590] <= r_data[18589];
                
                r_data[18591] <= r_data[18590];
                
                r_data[18592] <= r_data[18591];
                
                r_data[18593] <= r_data[18592];
                
                r_data[18594] <= r_data[18593];
                
                r_data[18595] <= r_data[18594];
                
                r_data[18596] <= r_data[18595];
                
                r_data[18597] <= r_data[18596];
                
                r_data[18598] <= r_data[18597];
                
                r_data[18599] <= r_data[18598];
                
                r_data[18600] <= r_data[18599];
                
                r_data[18601] <= r_data[18600];
                
                r_data[18602] <= r_data[18601];
                
                r_data[18603] <= r_data[18602];
                
                r_data[18604] <= r_data[18603];
                
                r_data[18605] <= r_data[18604];
                
                r_data[18606] <= r_data[18605];
                
                r_data[18607] <= r_data[18606];
                
                r_data[18608] <= r_data[18607];
                
                r_data[18609] <= r_data[18608];
                
                r_data[18610] <= r_data[18609];
                
                r_data[18611] <= r_data[18610];
                
                r_data[18612] <= r_data[18611];
                
                r_data[18613] <= r_data[18612];
                
                r_data[18614] <= r_data[18613];
                
                r_data[18615] <= r_data[18614];
                
                r_data[18616] <= r_data[18615];
                
                r_data[18617] <= r_data[18616];
                
                r_data[18618] <= r_data[18617];
                
                r_data[18619] <= r_data[18618];
                
                r_data[18620] <= r_data[18619];
                
                r_data[18621] <= r_data[18620];
                
                r_data[18622] <= r_data[18621];
                
                r_data[18623] <= r_data[18622];
                
                r_data[18624] <= r_data[18623];
                
                r_data[18625] <= r_data[18624];
                
                r_data[18626] <= r_data[18625];
                
                r_data[18627] <= r_data[18626];
                
                r_data[18628] <= r_data[18627];
                
                r_data[18629] <= r_data[18628];
                
                r_data[18630] <= r_data[18629];
                
                r_data[18631] <= r_data[18630];
                
                r_data[18632] <= r_data[18631];
                
                r_data[18633] <= r_data[18632];
                
                r_data[18634] <= r_data[18633];
                
                r_data[18635] <= r_data[18634];
                
                r_data[18636] <= r_data[18635];
                
                r_data[18637] <= r_data[18636];
                
                r_data[18638] <= r_data[18637];
                
                r_data[18639] <= r_data[18638];
                
                r_data[18640] <= r_data[18639];
                
                r_data[18641] <= r_data[18640];
                
                r_data[18642] <= r_data[18641];
                
                r_data[18643] <= r_data[18642];
                
                r_data[18644] <= r_data[18643];
                
                r_data[18645] <= r_data[18644];
                
                r_data[18646] <= r_data[18645];
                
                r_data[18647] <= r_data[18646];
                
                r_data[18648] <= r_data[18647];
                
                r_data[18649] <= r_data[18648];
                
                r_data[18650] <= r_data[18649];
                
                r_data[18651] <= r_data[18650];
                
                r_data[18652] <= r_data[18651];
                
                r_data[18653] <= r_data[18652];
                
                r_data[18654] <= r_data[18653];
                
                r_data[18655] <= r_data[18654];
                
                r_data[18656] <= r_data[18655];
                
                r_data[18657] <= r_data[18656];
                
                r_data[18658] <= r_data[18657];
                
                r_data[18659] <= r_data[18658];
                
                r_data[18660] <= r_data[18659];
                
                r_data[18661] <= r_data[18660];
                
                r_data[18662] <= r_data[18661];
                
                r_data[18663] <= r_data[18662];
                
                r_data[18664] <= r_data[18663];
                
                r_data[18665] <= r_data[18664];
                
                r_data[18666] <= r_data[18665];
                
                r_data[18667] <= r_data[18666];
                
                r_data[18668] <= r_data[18667];
                
                r_data[18669] <= r_data[18668];
                
                r_data[18670] <= r_data[18669];
                
                r_data[18671] <= r_data[18670];
                
                r_data[18672] <= r_data[18671];
                
                r_data[18673] <= r_data[18672];
                
                r_data[18674] <= r_data[18673];
                
                r_data[18675] <= r_data[18674];
                
                r_data[18676] <= r_data[18675];
                
                r_data[18677] <= r_data[18676];
                
                r_data[18678] <= r_data[18677];
                
                r_data[18679] <= r_data[18678];
                
                r_data[18680] <= r_data[18679];
                
                r_data[18681] <= r_data[18680];
                
                r_data[18682] <= r_data[18681];
                
                r_data[18683] <= r_data[18682];
                
                r_data[18684] <= r_data[18683];
                
                r_data[18685] <= r_data[18684];
                
                r_data[18686] <= r_data[18685];
                
                r_data[18687] <= r_data[18686];
                
                r_data[18688] <= r_data[18687];
                
                r_data[18689] <= r_data[18688];
                
                r_data[18690] <= r_data[18689];
                
                r_data[18691] <= r_data[18690];
                
                r_data[18692] <= r_data[18691];
                
                r_data[18693] <= r_data[18692];
                
                r_data[18694] <= r_data[18693];
                
                r_data[18695] <= r_data[18694];
                
                r_data[18696] <= r_data[18695];
                
                r_data[18697] <= r_data[18696];
                
                r_data[18698] <= r_data[18697];
                
                r_data[18699] <= r_data[18698];
                
                r_data[18700] <= r_data[18699];
                
                r_data[18701] <= r_data[18700];
                
                r_data[18702] <= r_data[18701];
                
                r_data[18703] <= r_data[18702];
                
                r_data[18704] <= r_data[18703];
                
                r_data[18705] <= r_data[18704];
                
                r_data[18706] <= r_data[18705];
                
                r_data[18707] <= r_data[18706];
                
                r_data[18708] <= r_data[18707];
                
                r_data[18709] <= r_data[18708];
                
                r_data[18710] <= r_data[18709];
                
                r_data[18711] <= r_data[18710];
                
                r_data[18712] <= r_data[18711];
                
                r_data[18713] <= r_data[18712];
                
                r_data[18714] <= r_data[18713];
                
                r_data[18715] <= r_data[18714];
                
                r_data[18716] <= r_data[18715];
                
                r_data[18717] <= r_data[18716];
                
                r_data[18718] <= r_data[18717];
                
                r_data[18719] <= r_data[18718];
                
                r_data[18720] <= r_data[18719];
                
                r_data[18721] <= r_data[18720];
                
                r_data[18722] <= r_data[18721];
                
                r_data[18723] <= r_data[18722];
                
                r_data[18724] <= r_data[18723];
                
                r_data[18725] <= r_data[18724];
                
                r_data[18726] <= r_data[18725];
                
                r_data[18727] <= r_data[18726];
                
                r_data[18728] <= r_data[18727];
                
                r_data[18729] <= r_data[18728];
                
                r_data[18730] <= r_data[18729];
                
                r_data[18731] <= r_data[18730];
                
                r_data[18732] <= r_data[18731];
                
                r_data[18733] <= r_data[18732];
                
                r_data[18734] <= r_data[18733];
                
                r_data[18735] <= r_data[18734];
                
                r_data[18736] <= r_data[18735];
                
                r_data[18737] <= r_data[18736];
                
                r_data[18738] <= r_data[18737];
                
                r_data[18739] <= r_data[18738];
                
                r_data[18740] <= r_data[18739];
                
                r_data[18741] <= r_data[18740];
                
                r_data[18742] <= r_data[18741];
                
                r_data[18743] <= r_data[18742];
                
                r_data[18744] <= r_data[18743];
                
                r_data[18745] <= r_data[18744];
                
                r_data[18746] <= r_data[18745];
                
                r_data[18747] <= r_data[18746];
                
                r_data[18748] <= r_data[18747];
                
                r_data[18749] <= r_data[18748];
                
                r_data[18750] <= r_data[18749];
                
                r_data[18751] <= r_data[18750];
                
                r_data[18752] <= r_data[18751];
                
                r_data[18753] <= r_data[18752];
                
                r_data[18754] <= r_data[18753];
                
                r_data[18755] <= r_data[18754];
                
                r_data[18756] <= r_data[18755];
                
                r_data[18757] <= r_data[18756];
                
                r_data[18758] <= r_data[18757];
                
                r_data[18759] <= r_data[18758];
                
                r_data[18760] <= r_data[18759];
                
                r_data[18761] <= r_data[18760];
                
                r_data[18762] <= r_data[18761];
                
                r_data[18763] <= r_data[18762];
                
                r_data[18764] <= r_data[18763];
                
                r_data[18765] <= r_data[18764];
                
                r_data[18766] <= r_data[18765];
                
                r_data[18767] <= r_data[18766];
                
                r_data[18768] <= r_data[18767];
                
                r_data[18769] <= r_data[18768];
                
                r_data[18770] <= r_data[18769];
                
                r_data[18771] <= r_data[18770];
                
                r_data[18772] <= r_data[18771];
                
                r_data[18773] <= r_data[18772];
                
                r_data[18774] <= r_data[18773];
                
                r_data[18775] <= r_data[18774];
                
                r_data[18776] <= r_data[18775];
                
                r_data[18777] <= r_data[18776];
                
                r_data[18778] <= r_data[18777];
                
                r_data[18779] <= r_data[18778];
                
                r_data[18780] <= r_data[18779];
                
                r_data[18781] <= r_data[18780];
                
                r_data[18782] <= r_data[18781];
                
                r_data[18783] <= r_data[18782];
                
                r_data[18784] <= r_data[18783];
                
                r_data[18785] <= r_data[18784];
                
                r_data[18786] <= r_data[18785];
                
                r_data[18787] <= r_data[18786];
                
                r_data[18788] <= r_data[18787];
                
                r_data[18789] <= r_data[18788];
                
                r_data[18790] <= r_data[18789];
                
                r_data[18791] <= r_data[18790];
                
                r_data[18792] <= r_data[18791];
                
                r_data[18793] <= r_data[18792];
                
                r_data[18794] <= r_data[18793];
                
                r_data[18795] <= r_data[18794];
                
                r_data[18796] <= r_data[18795];
                
                r_data[18797] <= r_data[18796];
                
                r_data[18798] <= r_data[18797];
                
                r_data[18799] <= r_data[18798];
                
                r_data[18800] <= r_data[18799];
                
                r_data[18801] <= r_data[18800];
                
                r_data[18802] <= r_data[18801];
                
                r_data[18803] <= r_data[18802];
                
                r_data[18804] <= r_data[18803];
                
                r_data[18805] <= r_data[18804];
                
                r_data[18806] <= r_data[18805];
                
                r_data[18807] <= r_data[18806];
                
                r_data[18808] <= r_data[18807];
                
                r_data[18809] <= r_data[18808];
                
                r_data[18810] <= r_data[18809];
                
                r_data[18811] <= r_data[18810];
                
                r_data[18812] <= r_data[18811];
                
                r_data[18813] <= r_data[18812];
                
                r_data[18814] <= r_data[18813];
                
                r_data[18815] <= r_data[18814];
                
                r_data[18816] <= r_data[18815];
                
                r_data[18817] <= r_data[18816];
                
                r_data[18818] <= r_data[18817];
                
                r_data[18819] <= r_data[18818];
                
                r_data[18820] <= r_data[18819];
                
                r_data[18821] <= r_data[18820];
                
                r_data[18822] <= r_data[18821];
                
                r_data[18823] <= r_data[18822];
                
                r_data[18824] <= r_data[18823];
                
                r_data[18825] <= r_data[18824];
                
                r_data[18826] <= r_data[18825];
                
                r_data[18827] <= r_data[18826];
                
                r_data[18828] <= r_data[18827];
                
                r_data[18829] <= r_data[18828];
                
                r_data[18830] <= r_data[18829];
                
                r_data[18831] <= r_data[18830];
                
                r_data[18832] <= r_data[18831];
                
                r_data[18833] <= r_data[18832];
                
                r_data[18834] <= r_data[18833];
                
                r_data[18835] <= r_data[18834];
                
                r_data[18836] <= r_data[18835];
                
                r_data[18837] <= r_data[18836];
                
                r_data[18838] <= r_data[18837];
                
                r_data[18839] <= r_data[18838];
                
                r_data[18840] <= r_data[18839];
                
                r_data[18841] <= r_data[18840];
                
                r_data[18842] <= r_data[18841];
                
                r_data[18843] <= r_data[18842];
                
                r_data[18844] <= r_data[18843];
                
                r_data[18845] <= r_data[18844];
                
                r_data[18846] <= r_data[18845];
                
                r_data[18847] <= r_data[18846];
                
                r_data[18848] <= r_data[18847];
                
                r_data[18849] <= r_data[18848];
                
                r_data[18850] <= r_data[18849];
                
                r_data[18851] <= r_data[18850];
                
                r_data[18852] <= r_data[18851];
                
                r_data[18853] <= r_data[18852];
                
                r_data[18854] <= r_data[18853];
                
                r_data[18855] <= r_data[18854];
                
                r_data[18856] <= r_data[18855];
                
                r_data[18857] <= r_data[18856];
                
                r_data[18858] <= r_data[18857];
                
                r_data[18859] <= r_data[18858];
                
                r_data[18860] <= r_data[18859];
                
                r_data[18861] <= r_data[18860];
                
                r_data[18862] <= r_data[18861];
                
                r_data[18863] <= r_data[18862];
                
                r_data[18864] <= r_data[18863];
                
                r_data[18865] <= r_data[18864];
                
                r_data[18866] <= r_data[18865];
                
                r_data[18867] <= r_data[18866];
                
                r_data[18868] <= r_data[18867];
                
                r_data[18869] <= r_data[18868];
                
                r_data[18870] <= r_data[18869];
                
                r_data[18871] <= r_data[18870];
                
                r_data[18872] <= r_data[18871];
                
                r_data[18873] <= r_data[18872];
                
                r_data[18874] <= r_data[18873];
                
                r_data[18875] <= r_data[18874];
                
                r_data[18876] <= r_data[18875];
                
                r_data[18877] <= r_data[18876];
                
                r_data[18878] <= r_data[18877];
                
                r_data[18879] <= r_data[18878];
                
                r_data[18880] <= r_data[18879];
                
                r_data[18881] <= r_data[18880];
                
                r_data[18882] <= r_data[18881];
                
                r_data[18883] <= r_data[18882];
                
                r_data[18884] <= r_data[18883];
                
                r_data[18885] <= r_data[18884];
                
                r_data[18886] <= r_data[18885];
                
                r_data[18887] <= r_data[18886];
                
                r_data[18888] <= r_data[18887];
                
                r_data[18889] <= r_data[18888];
                
                r_data[18890] <= r_data[18889];
                
                r_data[18891] <= r_data[18890];
                
                r_data[18892] <= r_data[18891];
                
                r_data[18893] <= r_data[18892];
                
                r_data[18894] <= r_data[18893];
                
                r_data[18895] <= r_data[18894];
                
                r_data[18896] <= r_data[18895];
                
                r_data[18897] <= r_data[18896];
                
                r_data[18898] <= r_data[18897];
                
                r_data[18899] <= r_data[18898];
                
                r_data[18900] <= r_data[18899];
                
                r_data[18901] <= r_data[18900];
                
                r_data[18902] <= r_data[18901];
                
                r_data[18903] <= r_data[18902];
                
                r_data[18904] <= r_data[18903];
                
                r_data[18905] <= r_data[18904];
                
                r_data[18906] <= r_data[18905];
                
                r_data[18907] <= r_data[18906];
                
                r_data[18908] <= r_data[18907];
                
                r_data[18909] <= r_data[18908];
                
                r_data[18910] <= r_data[18909];
                
                r_data[18911] <= r_data[18910];
                
                r_data[18912] <= r_data[18911];
                
                r_data[18913] <= r_data[18912];
                
                r_data[18914] <= r_data[18913];
                
                r_data[18915] <= r_data[18914];
                
                r_data[18916] <= r_data[18915];
                
                r_data[18917] <= r_data[18916];
                
                r_data[18918] <= r_data[18917];
                
                r_data[18919] <= r_data[18918];
                
                r_data[18920] <= r_data[18919];
                
                r_data[18921] <= r_data[18920];
                
                r_data[18922] <= r_data[18921];
                
                r_data[18923] <= r_data[18922];
                
                r_data[18924] <= r_data[18923];
                
                r_data[18925] <= r_data[18924];
                
                r_data[18926] <= r_data[18925];
                
                r_data[18927] <= r_data[18926];
                
                r_data[18928] <= r_data[18927];
                
                r_data[18929] <= r_data[18928];
                
                r_data[18930] <= r_data[18929];
                
                r_data[18931] <= r_data[18930];
                
                r_data[18932] <= r_data[18931];
                
                r_data[18933] <= r_data[18932];
                
                r_data[18934] <= r_data[18933];
                
                r_data[18935] <= r_data[18934];
                
                r_data[18936] <= r_data[18935];
                
                r_data[18937] <= r_data[18936];
                
                r_data[18938] <= r_data[18937];
                
                r_data[18939] <= r_data[18938];
                
                r_data[18940] <= r_data[18939];
                
                r_data[18941] <= r_data[18940];
                
                r_data[18942] <= r_data[18941];
                
                r_data[18943] <= r_data[18942];
                
                r_data[18944] <= r_data[18943];
                
                r_data[18945] <= r_data[18944];
                
                r_data[18946] <= r_data[18945];
                
                r_data[18947] <= r_data[18946];
                
                r_data[18948] <= r_data[18947];
                
                r_data[18949] <= r_data[18948];
                
                r_data[18950] <= r_data[18949];
                
                r_data[18951] <= r_data[18950];
                
                r_data[18952] <= r_data[18951];
                
                r_data[18953] <= r_data[18952];
                
                r_data[18954] <= r_data[18953];
                
                r_data[18955] <= r_data[18954];
                
                r_data[18956] <= r_data[18955];
                
                r_data[18957] <= r_data[18956];
                
                r_data[18958] <= r_data[18957];
                
                r_data[18959] <= r_data[18958];
                
                r_data[18960] <= r_data[18959];
                
                r_data[18961] <= r_data[18960];
                
                r_data[18962] <= r_data[18961];
                
                r_data[18963] <= r_data[18962];
                
                r_data[18964] <= r_data[18963];
                
                r_data[18965] <= r_data[18964];
                
                r_data[18966] <= r_data[18965];
                
                r_data[18967] <= r_data[18966];
                
                r_data[18968] <= r_data[18967];
                
                r_data[18969] <= r_data[18968];
                
                r_data[18970] <= r_data[18969];
                
                r_data[18971] <= r_data[18970];
                
                r_data[18972] <= r_data[18971];
                
                r_data[18973] <= r_data[18972];
                
                r_data[18974] <= r_data[18973];
                
                r_data[18975] <= r_data[18974];
                
                r_data[18976] <= r_data[18975];
                
                r_data[18977] <= r_data[18976];
                
                r_data[18978] <= r_data[18977];
                
                r_data[18979] <= r_data[18978];
                
                r_data[18980] <= r_data[18979];
                
                r_data[18981] <= r_data[18980];
                
                r_data[18982] <= r_data[18981];
                
                r_data[18983] <= r_data[18982];
                
                r_data[18984] <= r_data[18983];
                
                r_data[18985] <= r_data[18984];
                
                r_data[18986] <= r_data[18985];
                
                r_data[18987] <= r_data[18986];
                
                r_data[18988] <= r_data[18987];
                
                r_data[18989] <= r_data[18988];
                
                r_data[18990] <= r_data[18989];
                
                r_data[18991] <= r_data[18990];
                
                r_data[18992] <= r_data[18991];
                
                r_data[18993] <= r_data[18992];
                
                r_data[18994] <= r_data[18993];
                
                r_data[18995] <= r_data[18994];
                
                r_data[18996] <= r_data[18995];
                
                r_data[18997] <= r_data[18996];
                
                r_data[18998] <= r_data[18997];
                
                r_data[18999] <= r_data[18998];
                
                r_data[19000] <= r_data[18999];
                
                r_data[19001] <= r_data[19000];
                
                r_data[19002] <= r_data[19001];
                
                r_data[19003] <= r_data[19002];
                
                r_data[19004] <= r_data[19003];
                
                r_data[19005] <= r_data[19004];
                
                r_data[19006] <= r_data[19005];
                
                r_data[19007] <= r_data[19006];
                
                r_data[19008] <= r_data[19007];
                
                r_data[19009] <= r_data[19008];
                
                r_data[19010] <= r_data[19009];
                
                r_data[19011] <= r_data[19010];
                
                r_data[19012] <= r_data[19011];
                
                r_data[19013] <= r_data[19012];
                
                r_data[19014] <= r_data[19013];
                
                r_data[19015] <= r_data[19014];
                
                r_data[19016] <= r_data[19015];
                
                r_data[19017] <= r_data[19016];
                
                r_data[19018] <= r_data[19017];
                
                r_data[19019] <= r_data[19018];
                
                r_data[19020] <= r_data[19019];
                
                r_data[19021] <= r_data[19020];
                
                r_data[19022] <= r_data[19021];
                
                r_data[19023] <= r_data[19022];
                
                r_data[19024] <= r_data[19023];
                
                r_data[19025] <= r_data[19024];
                
                r_data[19026] <= r_data[19025];
                
                r_data[19027] <= r_data[19026];
                
                r_data[19028] <= r_data[19027];
                
                r_data[19029] <= r_data[19028];
                
                r_data[19030] <= r_data[19029];
                
                r_data[19031] <= r_data[19030];
                
                r_data[19032] <= r_data[19031];
                
                r_data[19033] <= r_data[19032];
                
                r_data[19034] <= r_data[19033];
                
                r_data[19035] <= r_data[19034];
                
                r_data[19036] <= r_data[19035];
                
                r_data[19037] <= r_data[19036];
                
                r_data[19038] <= r_data[19037];
                
                r_data[19039] <= r_data[19038];
                
                r_data[19040] <= r_data[19039];
                
                r_data[19041] <= r_data[19040];
                
                r_data[19042] <= r_data[19041];
                
                r_data[19043] <= r_data[19042];
                
                r_data[19044] <= r_data[19043];
                
                r_data[19045] <= r_data[19044];
                
                r_data[19046] <= r_data[19045];
                
                r_data[19047] <= r_data[19046];
                
                r_data[19048] <= r_data[19047];
                
                r_data[19049] <= r_data[19048];
                
                r_data[19050] <= r_data[19049];
                
                r_data[19051] <= r_data[19050];
                
                r_data[19052] <= r_data[19051];
                
                r_data[19053] <= r_data[19052];
                
                r_data[19054] <= r_data[19053];
                
                r_data[19055] <= r_data[19054];
                
                r_data[19056] <= r_data[19055];
                
                r_data[19057] <= r_data[19056];
                
                r_data[19058] <= r_data[19057];
                
                r_data[19059] <= r_data[19058];
                
                r_data[19060] <= r_data[19059];
                
                r_data[19061] <= r_data[19060];
                
                r_data[19062] <= r_data[19061];
                
                r_data[19063] <= r_data[19062];
                
                r_data[19064] <= r_data[19063];
                
                r_data[19065] <= r_data[19064];
                
                r_data[19066] <= r_data[19065];
                
                r_data[19067] <= r_data[19066];
                
                r_data[19068] <= r_data[19067];
                
                r_data[19069] <= r_data[19068];
                
                r_data[19070] <= r_data[19069];
                
                r_data[19071] <= r_data[19070];
                
                r_data[19072] <= r_data[19071];
                
                r_data[19073] <= r_data[19072];
                
                r_data[19074] <= r_data[19073];
                
                r_data[19075] <= r_data[19074];
                
                r_data[19076] <= r_data[19075];
                
                r_data[19077] <= r_data[19076];
                
                r_data[19078] <= r_data[19077];
                
                r_data[19079] <= r_data[19078];
                
                r_data[19080] <= r_data[19079];
                
                r_data[19081] <= r_data[19080];
                
                r_data[19082] <= r_data[19081];
                
                r_data[19083] <= r_data[19082];
                
                r_data[19084] <= r_data[19083];
                
                r_data[19085] <= r_data[19084];
                
                r_data[19086] <= r_data[19085];
                
                r_data[19087] <= r_data[19086];
                
                r_data[19088] <= r_data[19087];
                
                r_data[19089] <= r_data[19088];
                
                r_data[19090] <= r_data[19089];
                
                r_data[19091] <= r_data[19090];
                
                r_data[19092] <= r_data[19091];
                
                r_data[19093] <= r_data[19092];
                
                r_data[19094] <= r_data[19093];
                
                r_data[19095] <= r_data[19094];
                
                r_data[19096] <= r_data[19095];
                
                r_data[19097] <= r_data[19096];
                
                r_data[19098] <= r_data[19097];
                
                r_data[19099] <= r_data[19098];
                
                r_data[19100] <= r_data[19099];
                
                r_data[19101] <= r_data[19100];
                
                r_data[19102] <= r_data[19101];
                
                r_data[19103] <= r_data[19102];
                
                r_data[19104] <= r_data[19103];
                
                r_data[19105] <= r_data[19104];
                
                r_data[19106] <= r_data[19105];
                
                r_data[19107] <= r_data[19106];
                
                r_data[19108] <= r_data[19107];
                
                r_data[19109] <= r_data[19108];
                
                r_data[19110] <= r_data[19109];
                
                r_data[19111] <= r_data[19110];
                
                r_data[19112] <= r_data[19111];
                
                r_data[19113] <= r_data[19112];
                
                r_data[19114] <= r_data[19113];
                
                r_data[19115] <= r_data[19114];
                
                r_data[19116] <= r_data[19115];
                
                r_data[19117] <= r_data[19116];
                
                r_data[19118] <= r_data[19117];
                
                r_data[19119] <= r_data[19118];
                
                r_data[19120] <= r_data[19119];
                
                r_data[19121] <= r_data[19120];
                
                r_data[19122] <= r_data[19121];
                
                r_data[19123] <= r_data[19122];
                
                r_data[19124] <= r_data[19123];
                
                r_data[19125] <= r_data[19124];
                
                r_data[19126] <= r_data[19125];
                
                r_data[19127] <= r_data[19126];
                
                r_data[19128] <= r_data[19127];
                
                r_data[19129] <= r_data[19128];
                
                r_data[19130] <= r_data[19129];
                
                r_data[19131] <= r_data[19130];
                
                r_data[19132] <= r_data[19131];
                
                r_data[19133] <= r_data[19132];
                
                r_data[19134] <= r_data[19133];
                
                r_data[19135] <= r_data[19134];
                
                r_data[19136] <= r_data[19135];
                
                r_data[19137] <= r_data[19136];
                
                r_data[19138] <= r_data[19137];
                
                r_data[19139] <= r_data[19138];
                
                r_data[19140] <= r_data[19139];
                
                r_data[19141] <= r_data[19140];
                
                r_data[19142] <= r_data[19141];
                
                r_data[19143] <= r_data[19142];
                
                r_data[19144] <= r_data[19143];
                
                r_data[19145] <= r_data[19144];
                
                r_data[19146] <= r_data[19145];
                
                r_data[19147] <= r_data[19146];
                
                r_data[19148] <= r_data[19147];
                
                r_data[19149] <= r_data[19148];
                
                r_data[19150] <= r_data[19149];
                
                r_data[19151] <= r_data[19150];
                
                r_data[19152] <= r_data[19151];
                
                r_data[19153] <= r_data[19152];
                
                r_data[19154] <= r_data[19153];
                
                r_data[19155] <= r_data[19154];
                
                r_data[19156] <= r_data[19155];
                
                r_data[19157] <= r_data[19156];
                
                r_data[19158] <= r_data[19157];
                
                r_data[19159] <= r_data[19158];
                
                r_data[19160] <= r_data[19159];
                
                r_data[19161] <= r_data[19160];
                
                r_data[19162] <= r_data[19161];
                
                r_data[19163] <= r_data[19162];
                
                r_data[19164] <= r_data[19163];
                
                r_data[19165] <= r_data[19164];
                
                r_data[19166] <= r_data[19165];
                
                r_data[19167] <= r_data[19166];
                
                r_data[19168] <= r_data[19167];
                
                r_data[19169] <= r_data[19168];
                
                r_data[19170] <= r_data[19169];
                
                r_data[19171] <= r_data[19170];
                
                r_data[19172] <= r_data[19171];
                
                r_data[19173] <= r_data[19172];
                
                r_data[19174] <= r_data[19173];
                
                r_data[19175] <= r_data[19174];
                
                r_data[19176] <= r_data[19175];
                
                r_data[19177] <= r_data[19176];
                
                r_data[19178] <= r_data[19177];
                
                r_data[19179] <= r_data[19178];
                
                r_data[19180] <= r_data[19179];
                
                r_data[19181] <= r_data[19180];
                
                r_data[19182] <= r_data[19181];
                
                r_data[19183] <= r_data[19182];
                
                r_data[19184] <= r_data[19183];
                
                r_data[19185] <= r_data[19184];
                
                r_data[19186] <= r_data[19185];
                
                r_data[19187] <= r_data[19186];
                
                r_data[19188] <= r_data[19187];
                
                r_data[19189] <= r_data[19188];
                
                r_data[19190] <= r_data[19189];
                
                r_data[19191] <= r_data[19190];
                
                r_data[19192] <= r_data[19191];
                
                r_data[19193] <= r_data[19192];
                
                r_data[19194] <= r_data[19193];
                
                r_data[19195] <= r_data[19194];
                
                r_data[19196] <= r_data[19195];
                
                r_data[19197] <= r_data[19196];
                
                r_data[19198] <= r_data[19197];
                
                r_data[19199] <= r_data[19198];
                
                r_data[19200] <= r_data[19199];
                
                r_data[19201] <= r_data[19200];
                
                r_data[19202] <= r_data[19201];
                
                r_data[19203] <= r_data[19202];
                
                r_data[19204] <= r_data[19203];
                
                r_data[19205] <= r_data[19204];
                
                r_data[19206] <= r_data[19205];
                
                r_data[19207] <= r_data[19206];
                
                r_data[19208] <= r_data[19207];
                
                r_data[19209] <= r_data[19208];
                
                r_data[19210] <= r_data[19209];
                
                r_data[19211] <= r_data[19210];
                
                r_data[19212] <= r_data[19211];
                
                r_data[19213] <= r_data[19212];
                
                r_data[19214] <= r_data[19213];
                
                r_data[19215] <= r_data[19214];
                
                r_data[19216] <= r_data[19215];
                
                r_data[19217] <= r_data[19216];
                
                r_data[19218] <= r_data[19217];
                
                r_data[19219] <= r_data[19218];
                
                r_data[19220] <= r_data[19219];
                
                r_data[19221] <= r_data[19220];
                
                r_data[19222] <= r_data[19221];
                
                r_data[19223] <= r_data[19222];
                
                r_data[19224] <= r_data[19223];
                
                r_data[19225] <= r_data[19224];
                
                r_data[19226] <= r_data[19225];
                
                r_data[19227] <= r_data[19226];
                
                r_data[19228] <= r_data[19227];
                
                r_data[19229] <= r_data[19228];
                
                r_data[19230] <= r_data[19229];
                
                r_data[19231] <= r_data[19230];
                
                r_data[19232] <= r_data[19231];
                
                r_data[19233] <= r_data[19232];
                
                r_data[19234] <= r_data[19233];
                
                r_data[19235] <= r_data[19234];
                
                r_data[19236] <= r_data[19235];
                
                r_data[19237] <= r_data[19236];
                
                r_data[19238] <= r_data[19237];
                
                r_data[19239] <= r_data[19238];
                
                r_data[19240] <= r_data[19239];
                
                r_data[19241] <= r_data[19240];
                
                r_data[19242] <= r_data[19241];
                
                r_data[19243] <= r_data[19242];
                
                r_data[19244] <= r_data[19243];
                
                r_data[19245] <= r_data[19244];
                
                r_data[19246] <= r_data[19245];
                
                r_data[19247] <= r_data[19246];
                
                r_data[19248] <= r_data[19247];
                
                r_data[19249] <= r_data[19248];
                
                r_data[19250] <= r_data[19249];
                
                r_data[19251] <= r_data[19250];
                
                r_data[19252] <= r_data[19251];
                
                r_data[19253] <= r_data[19252];
                
                r_data[19254] <= r_data[19253];
                
                r_data[19255] <= r_data[19254];
                
                r_data[19256] <= r_data[19255];
                
                r_data[19257] <= r_data[19256];
                
                r_data[19258] <= r_data[19257];
                
                r_data[19259] <= r_data[19258];
                
                r_data[19260] <= r_data[19259];
                
                r_data[19261] <= r_data[19260];
                
                r_data[19262] <= r_data[19261];
                
                r_data[19263] <= r_data[19262];
                
                r_data[19264] <= r_data[19263];
                
                r_data[19265] <= r_data[19264];
                
                r_data[19266] <= r_data[19265];
                
                r_data[19267] <= r_data[19266];
                
                r_data[19268] <= r_data[19267];
                
                r_data[19269] <= r_data[19268];
                
                r_data[19270] <= r_data[19269];
                
                r_data[19271] <= r_data[19270];
                
                r_data[19272] <= r_data[19271];
                
                r_data[19273] <= r_data[19272];
                
                r_data[19274] <= r_data[19273];
                
                r_data[19275] <= r_data[19274];
                
                r_data[19276] <= r_data[19275];
                
                r_data[19277] <= r_data[19276];
                
                r_data[19278] <= r_data[19277];
                
                r_data[19279] <= r_data[19278];
                
                r_data[19280] <= r_data[19279];
                
                r_data[19281] <= r_data[19280];
                
                r_data[19282] <= r_data[19281];
                
                r_data[19283] <= r_data[19282];
                
                r_data[19284] <= r_data[19283];
                
                r_data[19285] <= r_data[19284];
                
                r_data[19286] <= r_data[19285];
                
                r_data[19287] <= r_data[19286];
                
                r_data[19288] <= r_data[19287];
                
                r_data[19289] <= r_data[19288];
                
                r_data[19290] <= r_data[19289];
                
                r_data[19291] <= r_data[19290];
                
                r_data[19292] <= r_data[19291];
                
                r_data[19293] <= r_data[19292];
                
                r_data[19294] <= r_data[19293];
                
                r_data[19295] <= r_data[19294];
                
                r_data[19296] <= r_data[19295];
                
                r_data[19297] <= r_data[19296];
                
                r_data[19298] <= r_data[19297];
                
                r_data[19299] <= r_data[19298];
                
                r_data[19300] <= r_data[19299];
                
                r_data[19301] <= r_data[19300];
                
                r_data[19302] <= r_data[19301];
                
                r_data[19303] <= r_data[19302];
                
                r_data[19304] <= r_data[19303];
                
                r_data[19305] <= r_data[19304];
                
                r_data[19306] <= r_data[19305];
                
                r_data[19307] <= r_data[19306];
                
                r_data[19308] <= r_data[19307];
                
                r_data[19309] <= r_data[19308];
                
                r_data[19310] <= r_data[19309];
                
                r_data[19311] <= r_data[19310];
                
                r_data[19312] <= r_data[19311];
                
                r_data[19313] <= r_data[19312];
                
                r_data[19314] <= r_data[19313];
                
                r_data[19315] <= r_data[19314];
                
                r_data[19316] <= r_data[19315];
                
                r_data[19317] <= r_data[19316];
                
                r_data[19318] <= r_data[19317];
                
                r_data[19319] <= r_data[19318];
                
                r_data[19320] <= r_data[19319];
                
                r_data[19321] <= r_data[19320];
                
                r_data[19322] <= r_data[19321];
                
                r_data[19323] <= r_data[19322];
                
                r_data[19324] <= r_data[19323];
                
                r_data[19325] <= r_data[19324];
                
                r_data[19326] <= r_data[19325];
                
                r_data[19327] <= r_data[19326];
                
                r_data[19328] <= r_data[19327];
                
                r_data[19329] <= r_data[19328];
                
                r_data[19330] <= r_data[19329];
                
                r_data[19331] <= r_data[19330];
                
                r_data[19332] <= r_data[19331];
                
                r_data[19333] <= r_data[19332];
                
                r_data[19334] <= r_data[19333];
                
                r_data[19335] <= r_data[19334];
                
                r_data[19336] <= r_data[19335];
                
                r_data[19337] <= r_data[19336];
                
                r_data[19338] <= r_data[19337];
                
                r_data[19339] <= r_data[19338];
                
                r_data[19340] <= r_data[19339];
                
                r_data[19341] <= r_data[19340];
                
                r_data[19342] <= r_data[19341];
                
                r_data[19343] <= r_data[19342];
                
                r_data[19344] <= r_data[19343];
                
                r_data[19345] <= r_data[19344];
                
                r_data[19346] <= r_data[19345];
                
                r_data[19347] <= r_data[19346];
                
                r_data[19348] <= r_data[19347];
                
                r_data[19349] <= r_data[19348];
                
                r_data[19350] <= r_data[19349];
                
                r_data[19351] <= r_data[19350];
                
                r_data[19352] <= r_data[19351];
                
                r_data[19353] <= r_data[19352];
                
                r_data[19354] <= r_data[19353];
                
                r_data[19355] <= r_data[19354];
                
                r_data[19356] <= r_data[19355];
                
                r_data[19357] <= r_data[19356];
                
                r_data[19358] <= r_data[19357];
                
                r_data[19359] <= r_data[19358];
                
                r_data[19360] <= r_data[19359];
                
                r_data[19361] <= r_data[19360];
                
                r_data[19362] <= r_data[19361];
                
                r_data[19363] <= r_data[19362];
                
                r_data[19364] <= r_data[19363];
                
                r_data[19365] <= r_data[19364];
                
                r_data[19366] <= r_data[19365];
                
                r_data[19367] <= r_data[19366];
                
                r_data[19368] <= r_data[19367];
                
                r_data[19369] <= r_data[19368];
                
                r_data[19370] <= r_data[19369];
                
                r_data[19371] <= r_data[19370];
                
                r_data[19372] <= r_data[19371];
                
                r_data[19373] <= r_data[19372];
                
                r_data[19374] <= r_data[19373];
                
                r_data[19375] <= r_data[19374];
                
                r_data[19376] <= r_data[19375];
                
                r_data[19377] <= r_data[19376];
                
                r_data[19378] <= r_data[19377];
                
                r_data[19379] <= r_data[19378];
                
                r_data[19380] <= r_data[19379];
                
                r_data[19381] <= r_data[19380];
                
                r_data[19382] <= r_data[19381];
                
                r_data[19383] <= r_data[19382];
                
                r_data[19384] <= r_data[19383];
                
                r_data[19385] <= r_data[19384];
                
                r_data[19386] <= r_data[19385];
                
                r_data[19387] <= r_data[19386];
                
                r_data[19388] <= r_data[19387];
                
                r_data[19389] <= r_data[19388];
                
                r_data[19390] <= r_data[19389];
                
                r_data[19391] <= r_data[19390];
                
                r_data[19392] <= r_data[19391];
                
                r_data[19393] <= r_data[19392];
                
                r_data[19394] <= r_data[19393];
                
                r_data[19395] <= r_data[19394];
                
                r_data[19396] <= r_data[19395];
                
                r_data[19397] <= r_data[19396];
                
                r_data[19398] <= r_data[19397];
                
                r_data[19399] <= r_data[19398];
                
                r_data[19400] <= r_data[19399];
                
                r_data[19401] <= r_data[19400];
                
                r_data[19402] <= r_data[19401];
                
                r_data[19403] <= r_data[19402];
                
                r_data[19404] <= r_data[19403];
                
                r_data[19405] <= r_data[19404];
                
                r_data[19406] <= r_data[19405];
                
                r_data[19407] <= r_data[19406];
                
                r_data[19408] <= r_data[19407];
                
                r_data[19409] <= r_data[19408];
                
                r_data[19410] <= r_data[19409];
                
                r_data[19411] <= r_data[19410];
                
                r_data[19412] <= r_data[19411];
                
                r_data[19413] <= r_data[19412];
                
                r_data[19414] <= r_data[19413];
                
                r_data[19415] <= r_data[19414];
                
                r_data[19416] <= r_data[19415];
                
                r_data[19417] <= r_data[19416];
                
                r_data[19418] <= r_data[19417];
                
                r_data[19419] <= r_data[19418];
                
                r_data[19420] <= r_data[19419];
                
                r_data[19421] <= r_data[19420];
                
                r_data[19422] <= r_data[19421];
                
                r_data[19423] <= r_data[19422];
                
                r_data[19424] <= r_data[19423];
                
                r_data[19425] <= r_data[19424];
                
                r_data[19426] <= r_data[19425];
                
                r_data[19427] <= r_data[19426];
                
                r_data[19428] <= r_data[19427];
                
                r_data[19429] <= r_data[19428];
                
                r_data[19430] <= r_data[19429];
                
                r_data[19431] <= r_data[19430];
                
                r_data[19432] <= r_data[19431];
                
                r_data[19433] <= r_data[19432];
                
                r_data[19434] <= r_data[19433];
                
                r_data[19435] <= r_data[19434];
                
                r_data[19436] <= r_data[19435];
                
                r_data[19437] <= r_data[19436];
                
                r_data[19438] <= r_data[19437];
                
                r_data[19439] <= r_data[19438];
                
                r_data[19440] <= r_data[19439];
                
                r_data[19441] <= r_data[19440];
                
                r_data[19442] <= r_data[19441];
                
                r_data[19443] <= r_data[19442];
                
                r_data[19444] <= r_data[19443];
                
                r_data[19445] <= r_data[19444];
                
                r_data[19446] <= r_data[19445];
                
                r_data[19447] <= r_data[19446];
                
                r_data[19448] <= r_data[19447];
                
                r_data[19449] <= r_data[19448];
                
                r_data[19450] <= r_data[19449];
                
                r_data[19451] <= r_data[19450];
                
                r_data[19452] <= r_data[19451];
                
                r_data[19453] <= r_data[19452];
                
                r_data[19454] <= r_data[19453];
                
                r_data[19455] <= r_data[19454];
                
                r_data[19456] <= r_data[19455];
                
                r_data[19457] <= r_data[19456];
                
                r_data[19458] <= r_data[19457];
                
                r_data[19459] <= r_data[19458];
                
                r_data[19460] <= r_data[19459];
                
                r_data[19461] <= r_data[19460];
                
                r_data[19462] <= r_data[19461];
                
                r_data[19463] <= r_data[19462];
                
                r_data[19464] <= r_data[19463];
                
                r_data[19465] <= r_data[19464];
                
                r_data[19466] <= r_data[19465];
                
                r_data[19467] <= r_data[19466];
                
                r_data[19468] <= r_data[19467];
                
                r_data[19469] <= r_data[19468];
                
                r_data[19470] <= r_data[19469];
                
                r_data[19471] <= r_data[19470];
                
                r_data[19472] <= r_data[19471];
                
                r_data[19473] <= r_data[19472];
                
                r_data[19474] <= r_data[19473];
                
                r_data[19475] <= r_data[19474];
                
                r_data[19476] <= r_data[19475];
                
                r_data[19477] <= r_data[19476];
                
                r_data[19478] <= r_data[19477];
                
                r_data[19479] <= r_data[19478];
                
                r_data[19480] <= r_data[19479];
                
                r_data[19481] <= r_data[19480];
                
                r_data[19482] <= r_data[19481];
                
                r_data[19483] <= r_data[19482];
                
                r_data[19484] <= r_data[19483];
                
                r_data[19485] <= r_data[19484];
                
                r_data[19486] <= r_data[19485];
                
                r_data[19487] <= r_data[19486];
                
                r_data[19488] <= r_data[19487];
                
                r_data[19489] <= r_data[19488];
                
                r_data[19490] <= r_data[19489];
                
                r_data[19491] <= r_data[19490];
                
                r_data[19492] <= r_data[19491];
                
                r_data[19493] <= r_data[19492];
                
                r_data[19494] <= r_data[19493];
                
                r_data[19495] <= r_data[19494];
                
                r_data[19496] <= r_data[19495];
                
                r_data[19497] <= r_data[19496];
                
                r_data[19498] <= r_data[19497];
                
                r_data[19499] <= r_data[19498];
                
                r_data[19500] <= r_data[19499];
                
                r_data[19501] <= r_data[19500];
                
                r_data[19502] <= r_data[19501];
                
                r_data[19503] <= r_data[19502];
                
                r_data[19504] <= r_data[19503];
                
                r_data[19505] <= r_data[19504];
                
                r_data[19506] <= r_data[19505];
                
                r_data[19507] <= r_data[19506];
                
                r_data[19508] <= r_data[19507];
                
                r_data[19509] <= r_data[19508];
                
                r_data[19510] <= r_data[19509];
                
                r_data[19511] <= r_data[19510];
                
                r_data[19512] <= r_data[19511];
                
                r_data[19513] <= r_data[19512];
                
                r_data[19514] <= r_data[19513];
                
                r_data[19515] <= r_data[19514];
                
                r_data[19516] <= r_data[19515];
                
                r_data[19517] <= r_data[19516];
                
                r_data[19518] <= r_data[19517];
                
                r_data[19519] <= r_data[19518];
                
                r_data[19520] <= r_data[19519];
                
                r_data[19521] <= r_data[19520];
                
                r_data[19522] <= r_data[19521];
                
                r_data[19523] <= r_data[19522];
                
                r_data[19524] <= r_data[19523];
                
                r_data[19525] <= r_data[19524];
                
                r_data[19526] <= r_data[19525];
                
                r_data[19527] <= r_data[19526];
                
                r_data[19528] <= r_data[19527];
                
                r_data[19529] <= r_data[19528];
                
                r_data[19530] <= r_data[19529];
                
                r_data[19531] <= r_data[19530];
                
                r_data[19532] <= r_data[19531];
                
                r_data[19533] <= r_data[19532];
                
                r_data[19534] <= r_data[19533];
                
                r_data[19535] <= r_data[19534];
                
                r_data[19536] <= r_data[19535];
                
                r_data[19537] <= r_data[19536];
                
                r_data[19538] <= r_data[19537];
                
                r_data[19539] <= r_data[19538];
                
                r_data[19540] <= r_data[19539];
                
                r_data[19541] <= r_data[19540];
                
                r_data[19542] <= r_data[19541];
                
                r_data[19543] <= r_data[19542];
                
                r_data[19544] <= r_data[19543];
                
                r_data[19545] <= r_data[19544];
                
                r_data[19546] <= r_data[19545];
                
                r_data[19547] <= r_data[19546];
                
                r_data[19548] <= r_data[19547];
                
                r_data[19549] <= r_data[19548];
                
                r_data[19550] <= r_data[19549];
                
                r_data[19551] <= r_data[19550];
                
                r_data[19552] <= r_data[19551];
                
                r_data[19553] <= r_data[19552];
                
                r_data[19554] <= r_data[19553];
                
                r_data[19555] <= r_data[19554];
                
                r_data[19556] <= r_data[19555];
                
                r_data[19557] <= r_data[19556];
                
                r_data[19558] <= r_data[19557];
                
                r_data[19559] <= r_data[19558];
                
                r_data[19560] <= r_data[19559];
                
                r_data[19561] <= r_data[19560];
                
                r_data[19562] <= r_data[19561];
                
                r_data[19563] <= r_data[19562];
                
                r_data[19564] <= r_data[19563];
                
                r_data[19565] <= r_data[19564];
                
                r_data[19566] <= r_data[19565];
                
                r_data[19567] <= r_data[19566];
                
                r_data[19568] <= r_data[19567];
                
                r_data[19569] <= r_data[19568];
                
                r_data[19570] <= r_data[19569];
                
                r_data[19571] <= r_data[19570];
                
                r_data[19572] <= r_data[19571];
                
                r_data[19573] <= r_data[19572];
                
                r_data[19574] <= r_data[19573];
                
                r_data[19575] <= r_data[19574];
                
                r_data[19576] <= r_data[19575];
                
                r_data[19577] <= r_data[19576];
                
                r_data[19578] <= r_data[19577];
                
                r_data[19579] <= r_data[19578];
                
                r_data[19580] <= r_data[19579];
                
                r_data[19581] <= r_data[19580];
                
                r_data[19582] <= r_data[19581];
                
                r_data[19583] <= r_data[19582];
                
                r_data[19584] <= r_data[19583];
                
                r_data[19585] <= r_data[19584];
                
                r_data[19586] <= r_data[19585];
                
                r_data[19587] <= r_data[19586];
                
                r_data[19588] <= r_data[19587];
                
                r_data[19589] <= r_data[19588];
                
                r_data[19590] <= r_data[19589];
                
                r_data[19591] <= r_data[19590];
                
                r_data[19592] <= r_data[19591];
                
                r_data[19593] <= r_data[19592];
                
                r_data[19594] <= r_data[19593];
                
                r_data[19595] <= r_data[19594];
                
                r_data[19596] <= r_data[19595];
                
                r_data[19597] <= r_data[19596];
                
                r_data[19598] <= r_data[19597];
                
                r_data[19599] <= r_data[19598];
                
                r_data[19600] <= r_data[19599];
                
                r_data[19601] <= r_data[19600];
                
                r_data[19602] <= r_data[19601];
                
                r_data[19603] <= r_data[19602];
                
                r_data[19604] <= r_data[19603];
                
                r_data[19605] <= r_data[19604];
                
                r_data[19606] <= r_data[19605];
                
                r_data[19607] <= r_data[19606];
                
                r_data[19608] <= r_data[19607];
                
                r_data[19609] <= r_data[19608];
                
                r_data[19610] <= r_data[19609];
                
                r_data[19611] <= r_data[19610];
                
                r_data[19612] <= r_data[19611];
                
                r_data[19613] <= r_data[19612];
                
                r_data[19614] <= r_data[19613];
                
                r_data[19615] <= r_data[19614];
                
                r_data[19616] <= r_data[19615];
                
                r_data[19617] <= r_data[19616];
                
                r_data[19618] <= r_data[19617];
                
                r_data[19619] <= r_data[19618];
                
                r_data[19620] <= r_data[19619];
                
                r_data[19621] <= r_data[19620];
                
                r_data[19622] <= r_data[19621];
                
                r_data[19623] <= r_data[19622];
                
                r_data[19624] <= r_data[19623];
                
                r_data[19625] <= r_data[19624];
                
                r_data[19626] <= r_data[19625];
                
                r_data[19627] <= r_data[19626];
                
                r_data[19628] <= r_data[19627];
                
                r_data[19629] <= r_data[19628];
                
                r_data[19630] <= r_data[19629];
                
                r_data[19631] <= r_data[19630];
                
                r_data[19632] <= r_data[19631];
                
                r_data[19633] <= r_data[19632];
                
                r_data[19634] <= r_data[19633];
                
                r_data[19635] <= r_data[19634];
                
                r_data[19636] <= r_data[19635];
                
                r_data[19637] <= r_data[19636];
                
                r_data[19638] <= r_data[19637];
                
                r_data[19639] <= r_data[19638];
                
                r_data[19640] <= r_data[19639];
                
                r_data[19641] <= r_data[19640];
                
                r_data[19642] <= r_data[19641];
                
                r_data[19643] <= r_data[19642];
                
                r_data[19644] <= r_data[19643];
                
                r_data[19645] <= r_data[19644];
                
                r_data[19646] <= r_data[19645];
                
                r_data[19647] <= r_data[19646];
                
                r_data[19648] <= r_data[19647];
                
                r_data[19649] <= r_data[19648];
                
                r_data[19650] <= r_data[19649];
                
                r_data[19651] <= r_data[19650];
                
                r_data[19652] <= r_data[19651];
                
                r_data[19653] <= r_data[19652];
                
                r_data[19654] <= r_data[19653];
                
                r_data[19655] <= r_data[19654];
                
                r_data[19656] <= r_data[19655];
                
                r_data[19657] <= r_data[19656];
                
                r_data[19658] <= r_data[19657];
                
                r_data[19659] <= r_data[19658];
                
                r_data[19660] <= r_data[19659];
                
                r_data[19661] <= r_data[19660];
                
                r_data[19662] <= r_data[19661];
                
                r_data[19663] <= r_data[19662];
                
                r_data[19664] <= r_data[19663];
                
                r_data[19665] <= r_data[19664];
                
                r_data[19666] <= r_data[19665];
                
                r_data[19667] <= r_data[19666];
                
                r_data[19668] <= r_data[19667];
                
                r_data[19669] <= r_data[19668];
                
                r_data[19670] <= r_data[19669];
                
                r_data[19671] <= r_data[19670];
                
                r_data[19672] <= r_data[19671];
                
                r_data[19673] <= r_data[19672];
                
                r_data[19674] <= r_data[19673];
                
                r_data[19675] <= r_data[19674];
                
                r_data[19676] <= r_data[19675];
                
                r_data[19677] <= r_data[19676];
                
                r_data[19678] <= r_data[19677];
                
                r_data[19679] <= r_data[19678];
                
                r_data[19680] <= r_data[19679];
                
                r_data[19681] <= r_data[19680];
                
                r_data[19682] <= r_data[19681];
                
                r_data[19683] <= r_data[19682];
                
                r_data[19684] <= r_data[19683];
                
                r_data[19685] <= r_data[19684];
                
                r_data[19686] <= r_data[19685];
                
                r_data[19687] <= r_data[19686];
                
                r_data[19688] <= r_data[19687];
                
                r_data[19689] <= r_data[19688];
                
                r_data[19690] <= r_data[19689];
                
                r_data[19691] <= r_data[19690];
                
                r_data[19692] <= r_data[19691];
                
                r_data[19693] <= r_data[19692];
                
                r_data[19694] <= r_data[19693];
                
                r_data[19695] <= r_data[19694];
                
                r_data[19696] <= r_data[19695];
                
                r_data[19697] <= r_data[19696];
                
                r_data[19698] <= r_data[19697];
                
                r_data[19699] <= r_data[19698];
                
                r_data[19700] <= r_data[19699];
                
                r_data[19701] <= r_data[19700];
                
                r_data[19702] <= r_data[19701];
                
                r_data[19703] <= r_data[19702];
                
                r_data[19704] <= r_data[19703];
                
                r_data[19705] <= r_data[19704];
                
                r_data[19706] <= r_data[19705];
                
                r_data[19707] <= r_data[19706];
                
                r_data[19708] <= r_data[19707];
                
                r_data[19709] <= r_data[19708];
                
                r_data[19710] <= r_data[19709];
                
                r_data[19711] <= r_data[19710];
                
                r_data[19712] <= r_data[19711];
                
                r_data[19713] <= r_data[19712];
                
                r_data[19714] <= r_data[19713];
                
                r_data[19715] <= r_data[19714];
                
                r_data[19716] <= r_data[19715];
                
                r_data[19717] <= r_data[19716];
                
                r_data[19718] <= r_data[19717];
                
                r_data[19719] <= r_data[19718];
                
                r_data[19720] <= r_data[19719];
                
                r_data[19721] <= r_data[19720];
                
                r_data[19722] <= r_data[19721];
                
                r_data[19723] <= r_data[19722];
                
                r_data[19724] <= r_data[19723];
                
                r_data[19725] <= r_data[19724];
                
                r_data[19726] <= r_data[19725];
                
                r_data[19727] <= r_data[19726];
                
                r_data[19728] <= r_data[19727];
                
                r_data[19729] <= r_data[19728];
                
                r_data[19730] <= r_data[19729];
                
                r_data[19731] <= r_data[19730];
                
                r_data[19732] <= r_data[19731];
                
                r_data[19733] <= r_data[19732];
                
                r_data[19734] <= r_data[19733];
                
                r_data[19735] <= r_data[19734];
                
                r_data[19736] <= r_data[19735];
                
                r_data[19737] <= r_data[19736];
                
                r_data[19738] <= r_data[19737];
                
                r_data[19739] <= r_data[19738];
                
                r_data[19740] <= r_data[19739];
                
                r_data[19741] <= r_data[19740];
                
                r_data[19742] <= r_data[19741];
                
                r_data[19743] <= r_data[19742];
                
                r_data[19744] <= r_data[19743];
                
                r_data[19745] <= r_data[19744];
                
                r_data[19746] <= r_data[19745];
                
                r_data[19747] <= r_data[19746];
                
                r_data[19748] <= r_data[19747];
                
                r_data[19749] <= r_data[19748];
                
                r_data[19750] <= r_data[19749];
                
                r_data[19751] <= r_data[19750];
                
                r_data[19752] <= r_data[19751];
                
                r_data[19753] <= r_data[19752];
                
                r_data[19754] <= r_data[19753];
                
                r_data[19755] <= r_data[19754];
                
                r_data[19756] <= r_data[19755];
                
                r_data[19757] <= r_data[19756];
                
                r_data[19758] <= r_data[19757];
                
                r_data[19759] <= r_data[19758];
                
                r_data[19760] <= r_data[19759];
                
                r_data[19761] <= r_data[19760];
                
                r_data[19762] <= r_data[19761];
                
                r_data[19763] <= r_data[19762];
                
                r_data[19764] <= r_data[19763];
                
                r_data[19765] <= r_data[19764];
                
                r_data[19766] <= r_data[19765];
                
                r_data[19767] <= r_data[19766];
                
                r_data[19768] <= r_data[19767];
                
                r_data[19769] <= r_data[19768];
                
                r_data[19770] <= r_data[19769];
                
                r_data[19771] <= r_data[19770];
                
                r_data[19772] <= r_data[19771];
                
                r_data[19773] <= r_data[19772];
                
                r_data[19774] <= r_data[19773];
                
                r_data[19775] <= r_data[19774];
                
                r_data[19776] <= r_data[19775];
                
                r_data[19777] <= r_data[19776];
                
                r_data[19778] <= r_data[19777];
                
                r_data[19779] <= r_data[19778];
                
                r_data[19780] <= r_data[19779];
                
                r_data[19781] <= r_data[19780];
                
                r_data[19782] <= r_data[19781];
                
                r_data[19783] <= r_data[19782];
                
                r_data[19784] <= r_data[19783];
                
                r_data[19785] <= r_data[19784];
                
                r_data[19786] <= r_data[19785];
                
                r_data[19787] <= r_data[19786];
                
                r_data[19788] <= r_data[19787];
                
                r_data[19789] <= r_data[19788];
                
                r_data[19790] <= r_data[19789];
                
                r_data[19791] <= r_data[19790];
                
                r_data[19792] <= r_data[19791];
                
                r_data[19793] <= r_data[19792];
                
                r_data[19794] <= r_data[19793];
                
                r_data[19795] <= r_data[19794];
                
                r_data[19796] <= r_data[19795];
                
                r_data[19797] <= r_data[19796];
                
                r_data[19798] <= r_data[19797];
                
                r_data[19799] <= r_data[19798];
                
                r_data[19800] <= r_data[19799];
                
                r_data[19801] <= r_data[19800];
                
                r_data[19802] <= r_data[19801];
                
                r_data[19803] <= r_data[19802];
                
                r_data[19804] <= r_data[19803];
                
                r_data[19805] <= r_data[19804];
                
                r_data[19806] <= r_data[19805];
                
                r_data[19807] <= r_data[19806];
                
                r_data[19808] <= r_data[19807];
                
                r_data[19809] <= r_data[19808];
                
                r_data[19810] <= r_data[19809];
                
                r_data[19811] <= r_data[19810];
                
                r_data[19812] <= r_data[19811];
                
                r_data[19813] <= r_data[19812];
                
                r_data[19814] <= r_data[19813];
                
                r_data[19815] <= r_data[19814];
                
                r_data[19816] <= r_data[19815];
                
                r_data[19817] <= r_data[19816];
                
                r_data[19818] <= r_data[19817];
                
                r_data[19819] <= r_data[19818];
                
                r_data[19820] <= r_data[19819];
                
                r_data[19821] <= r_data[19820];
                
                r_data[19822] <= r_data[19821];
                
                r_data[19823] <= r_data[19822];
                
                r_data[19824] <= r_data[19823];
                
                r_data[19825] <= r_data[19824];
                
                r_data[19826] <= r_data[19825];
                
                r_data[19827] <= r_data[19826];
                
                r_data[19828] <= r_data[19827];
                
                r_data[19829] <= r_data[19828];
                
                r_data[19830] <= r_data[19829];
                
                r_data[19831] <= r_data[19830];
                
                r_data[19832] <= r_data[19831];
                
                r_data[19833] <= r_data[19832];
                
                r_data[19834] <= r_data[19833];
                
                r_data[19835] <= r_data[19834];
                
                r_data[19836] <= r_data[19835];
                
                r_data[19837] <= r_data[19836];
                
                r_data[19838] <= r_data[19837];
                
                r_data[19839] <= r_data[19838];
                
                r_data[19840] <= r_data[19839];
                
                r_data[19841] <= r_data[19840];
                
                r_data[19842] <= r_data[19841];
                
                r_data[19843] <= r_data[19842];
                
                r_data[19844] <= r_data[19843];
                
                r_data[19845] <= r_data[19844];
                
                r_data[19846] <= r_data[19845];
                
                r_data[19847] <= r_data[19846];
                
                r_data[19848] <= r_data[19847];
                
                r_data[19849] <= r_data[19848];
                
                r_data[19850] <= r_data[19849];
                
                r_data[19851] <= r_data[19850];
                
                r_data[19852] <= r_data[19851];
                
                r_data[19853] <= r_data[19852];
                
                r_data[19854] <= r_data[19853];
                
                r_data[19855] <= r_data[19854];
                
                r_data[19856] <= r_data[19855];
                
                r_data[19857] <= r_data[19856];
                
                r_data[19858] <= r_data[19857];
                
                r_data[19859] <= r_data[19858];
                
                r_data[19860] <= r_data[19859];
                
                r_data[19861] <= r_data[19860];
                
                r_data[19862] <= r_data[19861];
                
                r_data[19863] <= r_data[19862];
                
                r_data[19864] <= r_data[19863];
                
                r_data[19865] <= r_data[19864];
                
                r_data[19866] <= r_data[19865];
                
                r_data[19867] <= r_data[19866];
                
                r_data[19868] <= r_data[19867];
                
                r_data[19869] <= r_data[19868];
                
                r_data[19870] <= r_data[19869];
                
                r_data[19871] <= r_data[19870];
                
                r_data[19872] <= r_data[19871];
                
                r_data[19873] <= r_data[19872];
                
                r_data[19874] <= r_data[19873];
                
                r_data[19875] <= r_data[19874];
                
                r_data[19876] <= r_data[19875];
                
                r_data[19877] <= r_data[19876];
                
                r_data[19878] <= r_data[19877];
                
                r_data[19879] <= r_data[19878];
                
                r_data[19880] <= r_data[19879];
                
                r_data[19881] <= r_data[19880];
                
                r_data[19882] <= r_data[19881];
                
                r_data[19883] <= r_data[19882];
                
                r_data[19884] <= r_data[19883];
                
                r_data[19885] <= r_data[19884];
                
                r_data[19886] <= r_data[19885];
                
                r_data[19887] <= r_data[19886];
                
                r_data[19888] <= r_data[19887];
                
                r_data[19889] <= r_data[19888];
                
                r_data[19890] <= r_data[19889];
                
                r_data[19891] <= r_data[19890];
                
                r_data[19892] <= r_data[19891];
                
                r_data[19893] <= r_data[19892];
                
                r_data[19894] <= r_data[19893];
                
                r_data[19895] <= r_data[19894];
                
                r_data[19896] <= r_data[19895];
                
                r_data[19897] <= r_data[19896];
                
                r_data[19898] <= r_data[19897];
                
                r_data[19899] <= r_data[19898];
                
                r_data[19900] <= r_data[19899];
                
                r_data[19901] <= r_data[19900];
                
                r_data[19902] <= r_data[19901];
                
                r_data[19903] <= r_data[19902];
                
                r_data[19904] <= r_data[19903];
                
                r_data[19905] <= r_data[19904];
                
                r_data[19906] <= r_data[19905];
                
                r_data[19907] <= r_data[19906];
                
                r_data[19908] <= r_data[19907];
                
                r_data[19909] <= r_data[19908];
                
                r_data[19910] <= r_data[19909];
                
                r_data[19911] <= r_data[19910];
                
                r_data[19912] <= r_data[19911];
                
                r_data[19913] <= r_data[19912];
                
                r_data[19914] <= r_data[19913];
                
                r_data[19915] <= r_data[19914];
                
                r_data[19916] <= r_data[19915];
                
                r_data[19917] <= r_data[19916];
                
                r_data[19918] <= r_data[19917];
                
                r_data[19919] <= r_data[19918];
                
                r_data[19920] <= r_data[19919];
                
                r_data[19921] <= r_data[19920];
                
                r_data[19922] <= r_data[19921];
                
                r_data[19923] <= r_data[19922];
                
                r_data[19924] <= r_data[19923];
                
                r_data[19925] <= r_data[19924];
                
                r_data[19926] <= r_data[19925];
                
                r_data[19927] <= r_data[19926];
                
                r_data[19928] <= r_data[19927];
                
                r_data[19929] <= r_data[19928];
                
                r_data[19930] <= r_data[19929];
                
                r_data[19931] <= r_data[19930];
                
                r_data[19932] <= r_data[19931];
                
                r_data[19933] <= r_data[19932];
                
                r_data[19934] <= r_data[19933];
                
                r_data[19935] <= r_data[19934];
                
                r_data[19936] <= r_data[19935];
                
                r_data[19937] <= r_data[19936];
                
                r_data[19938] <= r_data[19937];
                
                r_data[19939] <= r_data[19938];
                
                r_data[19940] <= r_data[19939];
                
                r_data[19941] <= r_data[19940];
                
                r_data[19942] <= r_data[19941];
                
                r_data[19943] <= r_data[19942];
                
                r_data[19944] <= r_data[19943];
                
                r_data[19945] <= r_data[19944];
                
                r_data[19946] <= r_data[19945];
                
                r_data[19947] <= r_data[19946];
                
                r_data[19948] <= r_data[19947];
                
                r_data[19949] <= r_data[19948];
                
                r_data[19950] <= r_data[19949];
                
                r_data[19951] <= r_data[19950];
                
                r_data[19952] <= r_data[19951];
                
                r_data[19953] <= r_data[19952];
                
                r_data[19954] <= r_data[19953];
                
                r_data[19955] <= r_data[19954];
                
                r_data[19956] <= r_data[19955];
                
                r_data[19957] <= r_data[19956];
                
                r_data[19958] <= r_data[19957];
                
                r_data[19959] <= r_data[19958];
                
                r_data[19960] <= r_data[19959];
                
                r_data[19961] <= r_data[19960];
                
                r_data[19962] <= r_data[19961];
                
                r_data[19963] <= r_data[19962];
                
                r_data[19964] <= r_data[19963];
                
                r_data[19965] <= r_data[19964];
                
                r_data[19966] <= r_data[19965];
                
                r_data[19967] <= r_data[19966];
                
                r_data[19968] <= r_data[19967];
                
                r_data[19969] <= r_data[19968];
                
                r_data[19970] <= r_data[19969];
                
                r_data[19971] <= r_data[19970];
                
                r_data[19972] <= r_data[19971];
                
                r_data[19973] <= r_data[19972];
                
                r_data[19974] <= r_data[19973];
                
                r_data[19975] <= r_data[19974];
                
                r_data[19976] <= r_data[19975];
                
                r_data[19977] <= r_data[19976];
                
                r_data[19978] <= r_data[19977];
                
                r_data[19979] <= r_data[19978];
                
                r_data[19980] <= r_data[19979];
                
                r_data[19981] <= r_data[19980];
                
                r_data[19982] <= r_data[19981];
                
                r_data[19983] <= r_data[19982];
                
                r_data[19984] <= r_data[19983];
                
                r_data[19985] <= r_data[19984];
                
                r_data[19986] <= r_data[19985];
                
                r_data[19987] <= r_data[19986];
                
                r_data[19988] <= r_data[19987];
                
                r_data[19989] <= r_data[19988];
                
                r_data[19990] <= r_data[19989];
                
                r_data[19991] <= r_data[19990];
                
                r_data[19992] <= r_data[19991];
                
                r_data[19993] <= r_data[19992];
                
                r_data[19994] <= r_data[19993];
                
                r_data[19995] <= r_data[19994];
                
                r_data[19996] <= r_data[19995];
                
                r_data[19997] <= r_data[19996];
                
                r_data[19998] <= r_data[19997];
                
                r_data[19999] <= r_data[19998];
                
                r_data[20000] <= r_data[19999];
                
                r_data[20001] <= r_data[20000];
                
                r_data[20002] <= r_data[20001];
                
                r_data[20003] <= r_data[20002];
                
                r_data[20004] <= r_data[20003];
                
                r_data[20005] <= r_data[20004];
                
                r_data[20006] <= r_data[20005];
                
                r_data[20007] <= r_data[20006];
                
                r_data[20008] <= r_data[20007];
                
                r_data[20009] <= r_data[20008];
                
                r_data[20010] <= r_data[20009];
                
                r_data[20011] <= r_data[20010];
                
                r_data[20012] <= r_data[20011];
                
                r_data[20013] <= r_data[20012];
                
                r_data[20014] <= r_data[20013];
                
                r_data[20015] <= r_data[20014];
                
                r_data[20016] <= r_data[20015];
                
                r_data[20017] <= r_data[20016];
                
                r_data[20018] <= r_data[20017];
                
                r_data[20019] <= r_data[20018];
                
                r_data[20020] <= r_data[20019];
                
                r_data[20021] <= r_data[20020];
                
                r_data[20022] <= r_data[20021];
                
                r_data[20023] <= r_data[20022];
                
                r_data[20024] <= r_data[20023];
                
                r_data[20025] <= r_data[20024];
                
                r_data[20026] <= r_data[20025];
                
                r_data[20027] <= r_data[20026];
                
                r_data[20028] <= r_data[20027];
                
                r_data[20029] <= r_data[20028];
                
                r_data[20030] <= r_data[20029];
                
                r_data[20031] <= r_data[20030];
                
                r_data[20032] <= r_data[20031];
                
                r_data[20033] <= r_data[20032];
                
                r_data[20034] <= r_data[20033];
                
                r_data[20035] <= r_data[20034];
                
                r_data[20036] <= r_data[20035];
                
                r_data[20037] <= r_data[20036];
                
                r_data[20038] <= r_data[20037];
                
                r_data[20039] <= r_data[20038];
                
                r_data[20040] <= r_data[20039];
                
                r_data[20041] <= r_data[20040];
                
                r_data[20042] <= r_data[20041];
                
                r_data[20043] <= r_data[20042];
                
                r_data[20044] <= r_data[20043];
                
                r_data[20045] <= r_data[20044];
                
                r_data[20046] <= r_data[20045];
                
                r_data[20047] <= r_data[20046];
                
                r_data[20048] <= r_data[20047];
                
                r_data[20049] <= r_data[20048];
                
                r_data[20050] <= r_data[20049];
                
                r_data[20051] <= r_data[20050];
                
                r_data[20052] <= r_data[20051];
                
                r_data[20053] <= r_data[20052];
                
                r_data[20054] <= r_data[20053];
                
                r_data[20055] <= r_data[20054];
                
                r_data[20056] <= r_data[20055];
                
                r_data[20057] <= r_data[20056];
                
                r_data[20058] <= r_data[20057];
                
                r_data[20059] <= r_data[20058];
                
                r_data[20060] <= r_data[20059];
                
                r_data[20061] <= r_data[20060];
                
                r_data[20062] <= r_data[20061];
                
                r_data[20063] <= r_data[20062];
                
                r_data[20064] <= r_data[20063];
                
                r_data[20065] <= r_data[20064];
                
                r_data[20066] <= r_data[20065];
                
                r_data[20067] <= r_data[20066];
                
                r_data[20068] <= r_data[20067];
                
                r_data[20069] <= r_data[20068];
                
                r_data[20070] <= r_data[20069];
                
                r_data[20071] <= r_data[20070];
                
                r_data[20072] <= r_data[20071];
                
                r_data[20073] <= r_data[20072];
                
                r_data[20074] <= r_data[20073];
                
                r_data[20075] <= r_data[20074];
                
                r_data[20076] <= r_data[20075];
                
                r_data[20077] <= r_data[20076];
                
                r_data[20078] <= r_data[20077];
                
                r_data[20079] <= r_data[20078];
                
                r_data[20080] <= r_data[20079];
                
                r_data[20081] <= r_data[20080];
                
                r_data[20082] <= r_data[20081];
                
                r_data[20083] <= r_data[20082];
                
                r_data[20084] <= r_data[20083];
                
                r_data[20085] <= r_data[20084];
                
                r_data[20086] <= r_data[20085];
                
                r_data[20087] <= r_data[20086];
                
                r_data[20088] <= r_data[20087];
                
                r_data[20089] <= r_data[20088];
                
                r_data[20090] <= r_data[20089];
                
                r_data[20091] <= r_data[20090];
                
                r_data[20092] <= r_data[20091];
                
                r_data[20093] <= r_data[20092];
                
                r_data[20094] <= r_data[20093];
                
                r_data[20095] <= r_data[20094];
                
                r_data[20096] <= r_data[20095];
                
                r_data[20097] <= r_data[20096];
                
                r_data[20098] <= r_data[20097];
                
                r_data[20099] <= r_data[20098];
                
                r_data[20100] <= r_data[20099];
                
                r_data[20101] <= r_data[20100];
                
                r_data[20102] <= r_data[20101];
                
                r_data[20103] <= r_data[20102];
                
                r_data[20104] <= r_data[20103];
                
                r_data[20105] <= r_data[20104];
                
                r_data[20106] <= r_data[20105];
                
                r_data[20107] <= r_data[20106];
                
                r_data[20108] <= r_data[20107];
                
                r_data[20109] <= r_data[20108];
                
                r_data[20110] <= r_data[20109];
                
                r_data[20111] <= r_data[20110];
                
                r_data[20112] <= r_data[20111];
                
                r_data[20113] <= r_data[20112];
                
                r_data[20114] <= r_data[20113];
                
                r_data[20115] <= r_data[20114];
                
                r_data[20116] <= r_data[20115];
                
                r_data[20117] <= r_data[20116];
                
                r_data[20118] <= r_data[20117];
                
                r_data[20119] <= r_data[20118];
                
                r_data[20120] <= r_data[20119];
                
                r_data[20121] <= r_data[20120];
                
                r_data[20122] <= r_data[20121];
                
                r_data[20123] <= r_data[20122];
                
                r_data[20124] <= r_data[20123];
                
                r_data[20125] <= r_data[20124];
                
                r_data[20126] <= r_data[20125];
                
                r_data[20127] <= r_data[20126];
                
                r_data[20128] <= r_data[20127];
                
                r_data[20129] <= r_data[20128];
                
                r_data[20130] <= r_data[20129];
                
                r_data[20131] <= r_data[20130];
                
                r_data[20132] <= r_data[20131];
                
                r_data[20133] <= r_data[20132];
                
                r_data[20134] <= r_data[20133];
                
                r_data[20135] <= r_data[20134];
                
                r_data[20136] <= r_data[20135];
                
                r_data[20137] <= r_data[20136];
                
                r_data[20138] <= r_data[20137];
                
                r_data[20139] <= r_data[20138];
                
                r_data[20140] <= r_data[20139];
                
                r_data[20141] <= r_data[20140];
                
                r_data[20142] <= r_data[20141];
                
                r_data[20143] <= r_data[20142];
                
                r_data[20144] <= r_data[20143];
                
                r_data[20145] <= r_data[20144];
                
                r_data[20146] <= r_data[20145];
                
                r_data[20147] <= r_data[20146];
                
                r_data[20148] <= r_data[20147];
                
                r_data[20149] <= r_data[20148];
                
                r_data[20150] <= r_data[20149];
                
                r_data[20151] <= r_data[20150];
                
                r_data[20152] <= r_data[20151];
                
                r_data[20153] <= r_data[20152];
                
                r_data[20154] <= r_data[20153];
                
                r_data[20155] <= r_data[20154];
                
                r_data[20156] <= r_data[20155];
                
                r_data[20157] <= r_data[20156];
                
                r_data[20158] <= r_data[20157];
                
                r_data[20159] <= r_data[20158];
                
                r_data[20160] <= r_data[20159];
                
                r_data[20161] <= r_data[20160];
                
                r_data[20162] <= r_data[20161];
                
                r_data[20163] <= r_data[20162];
                
                r_data[20164] <= r_data[20163];
                
                r_data[20165] <= r_data[20164];
                
                r_data[20166] <= r_data[20165];
                
                r_data[20167] <= r_data[20166];
                
                r_data[20168] <= r_data[20167];
                
                r_data[20169] <= r_data[20168];
                
                r_data[20170] <= r_data[20169];
                
                r_data[20171] <= r_data[20170];
                
                r_data[20172] <= r_data[20171];
                
                r_data[20173] <= r_data[20172];
                
                r_data[20174] <= r_data[20173];
                
                r_data[20175] <= r_data[20174];
                
                r_data[20176] <= r_data[20175];
                
                r_data[20177] <= r_data[20176];
                
                r_data[20178] <= r_data[20177];
                
                r_data[20179] <= r_data[20178];
                
                r_data[20180] <= r_data[20179];
                
                r_data[20181] <= r_data[20180];
                
                r_data[20182] <= r_data[20181];
                
                r_data[20183] <= r_data[20182];
                
                r_data[20184] <= r_data[20183];
                
                r_data[20185] <= r_data[20184];
                
                r_data[20186] <= r_data[20185];
                
                r_data[20187] <= r_data[20186];
                
                r_data[20188] <= r_data[20187];
                
                r_data[20189] <= r_data[20188];
                
                r_data[20190] <= r_data[20189];
                
                r_data[20191] <= r_data[20190];
                
                r_data[20192] <= r_data[20191];
                
                r_data[20193] <= r_data[20192];
                
                r_data[20194] <= r_data[20193];
                
                r_data[20195] <= r_data[20194];
                
                r_data[20196] <= r_data[20195];
                
                r_data[20197] <= r_data[20196];
                
                r_data[20198] <= r_data[20197];
                
                r_data[20199] <= r_data[20198];
                
                r_data[20200] <= r_data[20199];
                
                r_data[20201] <= r_data[20200];
                
                r_data[20202] <= r_data[20201];
                
                r_data[20203] <= r_data[20202];
                
                r_data[20204] <= r_data[20203];
                
                r_data[20205] <= r_data[20204];
                
                r_data[20206] <= r_data[20205];
                
                r_data[20207] <= r_data[20206];
                
                r_data[20208] <= r_data[20207];
                
                r_data[20209] <= r_data[20208];
                
                r_data[20210] <= r_data[20209];
                
                r_data[20211] <= r_data[20210];
                
                r_data[20212] <= r_data[20211];
                
                r_data[20213] <= r_data[20212];
                
                r_data[20214] <= r_data[20213];
                
                r_data[20215] <= r_data[20214];
                
                r_data[20216] <= r_data[20215];
                
                r_data[20217] <= r_data[20216];
                
                r_data[20218] <= r_data[20217];
                
                r_data[20219] <= r_data[20218];
                
                r_data[20220] <= r_data[20219];
                
                r_data[20221] <= r_data[20220];
                
                r_data[20222] <= r_data[20221];
                
                r_data[20223] <= r_data[20222];
                
                r_data[20224] <= r_data[20223];
                
                r_data[20225] <= r_data[20224];
                
                r_data[20226] <= r_data[20225];
                
                r_data[20227] <= r_data[20226];
                
                r_data[20228] <= r_data[20227];
                
                r_data[20229] <= r_data[20228];
                
                r_data[20230] <= r_data[20229];
                
                r_data[20231] <= r_data[20230];
                
                r_data[20232] <= r_data[20231];
                
                r_data[20233] <= r_data[20232];
                
                r_data[20234] <= r_data[20233];
                
                r_data[20235] <= r_data[20234];
                
                r_data[20236] <= r_data[20235];
                
                r_data[20237] <= r_data[20236];
                
                r_data[20238] <= r_data[20237];
                
                r_data[20239] <= r_data[20238];
                
                r_data[20240] <= r_data[20239];
                
                r_data[20241] <= r_data[20240];
                
                r_data[20242] <= r_data[20241];
                
                r_data[20243] <= r_data[20242];
                
                r_data[20244] <= r_data[20243];
                
                r_data[20245] <= r_data[20244];
                
                r_data[20246] <= r_data[20245];
                
                r_data[20247] <= r_data[20246];
                
                r_data[20248] <= r_data[20247];
                
                r_data[20249] <= r_data[20248];
                
                r_data[20250] <= r_data[20249];
                
                r_data[20251] <= r_data[20250];
                
                r_data[20252] <= r_data[20251];
                
                r_data[20253] <= r_data[20252];
                
                r_data[20254] <= r_data[20253];
                
                r_data[20255] <= r_data[20254];
                
                r_data[20256] <= r_data[20255];
                
                r_data[20257] <= r_data[20256];
                
                r_data[20258] <= r_data[20257];
                
                r_data[20259] <= r_data[20258];
                
                r_data[20260] <= r_data[20259];
                
                r_data[20261] <= r_data[20260];
                
                r_data[20262] <= r_data[20261];
                
                r_data[20263] <= r_data[20262];
                
                r_data[20264] <= r_data[20263];
                
                r_data[20265] <= r_data[20264];
                
                r_data[20266] <= r_data[20265];
                
                r_data[20267] <= r_data[20266];
                
                r_data[20268] <= r_data[20267];
                
                r_data[20269] <= r_data[20268];
                
                r_data[20270] <= r_data[20269];
                
                r_data[20271] <= r_data[20270];
                
                r_data[20272] <= r_data[20271];
                
                r_data[20273] <= r_data[20272];
                
                r_data[20274] <= r_data[20273];
                
                r_data[20275] <= r_data[20274];
                
                r_data[20276] <= r_data[20275];
                
                r_data[20277] <= r_data[20276];
                
                r_data[20278] <= r_data[20277];
                
                r_data[20279] <= r_data[20278];
                
                r_data[20280] <= r_data[20279];
                
                r_data[20281] <= r_data[20280];
                
                r_data[20282] <= r_data[20281];
                
                r_data[20283] <= r_data[20282];
                
                r_data[20284] <= r_data[20283];
                
                r_data[20285] <= r_data[20284];
                
                r_data[20286] <= r_data[20285];
                
                r_data[20287] <= r_data[20286];
                
                r_data[20288] <= r_data[20287];
                
                r_data[20289] <= r_data[20288];
                
                r_data[20290] <= r_data[20289];
                
                r_data[20291] <= r_data[20290];
                
                r_data[20292] <= r_data[20291];
                
                r_data[20293] <= r_data[20292];
                
                r_data[20294] <= r_data[20293];
                
                r_data[20295] <= r_data[20294];
                
                r_data[20296] <= r_data[20295];
                
                r_data[20297] <= r_data[20296];
                
                r_data[20298] <= r_data[20297];
                
                r_data[20299] <= r_data[20298];
                
                r_data[20300] <= r_data[20299];
                
                r_data[20301] <= r_data[20300];
                
                r_data[20302] <= r_data[20301];
                
                r_data[20303] <= r_data[20302];
                
                r_data[20304] <= r_data[20303];
                
                r_data[20305] <= r_data[20304];
                
                r_data[20306] <= r_data[20305];
                
                r_data[20307] <= r_data[20306];
                
                r_data[20308] <= r_data[20307];
                
                r_data[20309] <= r_data[20308];
                
                r_data[20310] <= r_data[20309];
                
                r_data[20311] <= r_data[20310];
                
                r_data[20312] <= r_data[20311];
                
                r_data[20313] <= r_data[20312];
                
                r_data[20314] <= r_data[20313];
                
                r_data[20315] <= r_data[20314];
                
                r_data[20316] <= r_data[20315];
                
                r_data[20317] <= r_data[20316];
                
                r_data[20318] <= r_data[20317];
                
                r_data[20319] <= r_data[20318];
                
                r_data[20320] <= r_data[20319];
                
                r_data[20321] <= r_data[20320];
                
                r_data[20322] <= r_data[20321];
                
                r_data[20323] <= r_data[20322];
                
                r_data[20324] <= r_data[20323];
                
                r_data[20325] <= r_data[20324];
                
                r_data[20326] <= r_data[20325];
                
                r_data[20327] <= r_data[20326];
                
                r_data[20328] <= r_data[20327];
                
                r_data[20329] <= r_data[20328];
                
                r_data[20330] <= r_data[20329];
                
                r_data[20331] <= r_data[20330];
                
                r_data[20332] <= r_data[20331];
                
                r_data[20333] <= r_data[20332];
                
                r_data[20334] <= r_data[20333];
                
                r_data[20335] <= r_data[20334];
                
                r_data[20336] <= r_data[20335];
                
                r_data[20337] <= r_data[20336];
                
                r_data[20338] <= r_data[20337];
                
                r_data[20339] <= r_data[20338];
                
                r_data[20340] <= r_data[20339];
                
                r_data[20341] <= r_data[20340];
                
                r_data[20342] <= r_data[20341];
                
                r_data[20343] <= r_data[20342];
                
                r_data[20344] <= r_data[20343];
                
                r_data[20345] <= r_data[20344];
                
                r_data[20346] <= r_data[20345];
                
                r_data[20347] <= r_data[20346];
                
                r_data[20348] <= r_data[20347];
                
                r_data[20349] <= r_data[20348];
                
                r_data[20350] <= r_data[20349];
                
                r_data[20351] <= r_data[20350];
                
                r_data[20352] <= r_data[20351];
                
                r_data[20353] <= r_data[20352];
                
                r_data[20354] <= r_data[20353];
                
                r_data[20355] <= r_data[20354];
                
                r_data[20356] <= r_data[20355];
                
                r_data[20357] <= r_data[20356];
                
                r_data[20358] <= r_data[20357];
                
                r_data[20359] <= r_data[20358];
                
                r_data[20360] <= r_data[20359];
                
                r_data[20361] <= r_data[20360];
                
                r_data[20362] <= r_data[20361];
                
                r_data[20363] <= r_data[20362];
                
                r_data[20364] <= r_data[20363];
                
                r_data[20365] <= r_data[20364];
                
                r_data[20366] <= r_data[20365];
                
                r_data[20367] <= r_data[20366];
                
                r_data[20368] <= r_data[20367];
                
                r_data[20369] <= r_data[20368];
                
                r_data[20370] <= r_data[20369];
                
                r_data[20371] <= r_data[20370];
                
                r_data[20372] <= r_data[20371];
                
                r_data[20373] <= r_data[20372];
                
                r_data[20374] <= r_data[20373];
                
                r_data[20375] <= r_data[20374];
                
                r_data[20376] <= r_data[20375];
                
                r_data[20377] <= r_data[20376];
                
                r_data[20378] <= r_data[20377];
                
                r_data[20379] <= r_data[20378];
                
                r_data[20380] <= r_data[20379];
                
                r_data[20381] <= r_data[20380];
                
                r_data[20382] <= r_data[20381];
                
                r_data[20383] <= r_data[20382];
                
                r_data[20384] <= r_data[20383];
                
                r_data[20385] <= r_data[20384];
                
                r_data[20386] <= r_data[20385];
                
                r_data[20387] <= r_data[20386];
                
                r_data[20388] <= r_data[20387];
                
                r_data[20389] <= r_data[20388];
                
                r_data[20390] <= r_data[20389];
                
                r_data[20391] <= r_data[20390];
                
                r_data[20392] <= r_data[20391];
                
                r_data[20393] <= r_data[20392];
                
                r_data[20394] <= r_data[20393];
                
                r_data[20395] <= r_data[20394];
                
                r_data[20396] <= r_data[20395];
                
                r_data[20397] <= r_data[20396];
                
                r_data[20398] <= r_data[20397];
                
                r_data[20399] <= r_data[20398];
                
                r_data[20400] <= r_data[20399];
                
                r_data[20401] <= r_data[20400];
                
                r_data[20402] <= r_data[20401];
                
                r_data[20403] <= r_data[20402];
                
                r_data[20404] <= r_data[20403];
                
                r_data[20405] <= r_data[20404];
                
                r_data[20406] <= r_data[20405];
                
                r_data[20407] <= r_data[20406];
                
                r_data[20408] <= r_data[20407];
                
                r_data[20409] <= r_data[20408];
                
                r_data[20410] <= r_data[20409];
                
                r_data[20411] <= r_data[20410];
                
                r_data[20412] <= r_data[20411];
                
                r_data[20413] <= r_data[20412];
                
                r_data[20414] <= r_data[20413];
                
                r_data[20415] <= r_data[20414];
                
                r_data[20416] <= r_data[20415];
                
                r_data[20417] <= r_data[20416];
                
                r_data[20418] <= r_data[20417];
                
                r_data[20419] <= r_data[20418];
                
                r_data[20420] <= r_data[20419];
                
                r_data[20421] <= r_data[20420];
                
                r_data[20422] <= r_data[20421];
                
                r_data[20423] <= r_data[20422];
                
                r_data[20424] <= r_data[20423];
                
                r_data[20425] <= r_data[20424];
                
                r_data[20426] <= r_data[20425];
                
                r_data[20427] <= r_data[20426];
                
                r_data[20428] <= r_data[20427];
                
                r_data[20429] <= r_data[20428];
                
                r_data[20430] <= r_data[20429];
                
                r_data[20431] <= r_data[20430];
                
                r_data[20432] <= r_data[20431];
                
                r_data[20433] <= r_data[20432];
                
                r_data[20434] <= r_data[20433];
                
                r_data[20435] <= r_data[20434];
                
                r_data[20436] <= r_data[20435];
                
                r_data[20437] <= r_data[20436];
                
                r_data[20438] <= r_data[20437];
                
                r_data[20439] <= r_data[20438];
                
                r_data[20440] <= r_data[20439];
                
                r_data[20441] <= r_data[20440];
                
                r_data[20442] <= r_data[20441];
                
                r_data[20443] <= r_data[20442];
                
                r_data[20444] <= r_data[20443];
                
                r_data[20445] <= r_data[20444];
                
                r_data[20446] <= r_data[20445];
                
                r_data[20447] <= r_data[20446];
                
                r_data[20448] <= r_data[20447];
                
                r_data[20449] <= r_data[20448];
                
                r_data[20450] <= r_data[20449];
                
                r_data[20451] <= r_data[20450];
                
                r_data[20452] <= r_data[20451];
                
                r_data[20453] <= r_data[20452];
                
                r_data[20454] <= r_data[20453];
                
                r_data[20455] <= r_data[20454];
                
                r_data[20456] <= r_data[20455];
                
                r_data[20457] <= r_data[20456];
                
                r_data[20458] <= r_data[20457];
                
                r_data[20459] <= r_data[20458];
                
                r_data[20460] <= r_data[20459];
                
                r_data[20461] <= r_data[20460];
                
                r_data[20462] <= r_data[20461];
                
                r_data[20463] <= r_data[20462];
                
                r_data[20464] <= r_data[20463];
                
                r_data[20465] <= r_data[20464];
                
                r_data[20466] <= r_data[20465];
                
                r_data[20467] <= r_data[20466];
                
                r_data[20468] <= r_data[20467];
                
                r_data[20469] <= r_data[20468];
                
                r_data[20470] <= r_data[20469];
                
                r_data[20471] <= r_data[20470];
                
                r_data[20472] <= r_data[20471];
                
                r_data[20473] <= r_data[20472];
                
                r_data[20474] <= r_data[20473];
                
                r_data[20475] <= r_data[20474];
                
                r_data[20476] <= r_data[20475];
                
                r_data[20477] <= r_data[20476];
                
                r_data[20478] <= r_data[20477];
                
                r_data[20479] <= r_data[20478];
                
                r_data[20480] <= r_data[20479];
                
                r_data[20481] <= r_data[20480];
                
                r_data[20482] <= r_data[20481];
                
                r_data[20483] <= r_data[20482];
                
                r_data[20484] <= r_data[20483];
                
                r_data[20485] <= r_data[20484];
                
                r_data[20486] <= r_data[20485];
                
                r_data[20487] <= r_data[20486];
                
                r_data[20488] <= r_data[20487];
                
                r_data[20489] <= r_data[20488];
                
                r_data[20490] <= r_data[20489];
                
                r_data[20491] <= r_data[20490];
                
                r_data[20492] <= r_data[20491];
                
                r_data[20493] <= r_data[20492];
                
                r_data[20494] <= r_data[20493];
                
                r_data[20495] <= r_data[20494];
                
                r_data[20496] <= r_data[20495];
                
                r_data[20497] <= r_data[20496];
                
                r_data[20498] <= r_data[20497];
                
                r_data[20499] <= r_data[20498];
                
                r_data[20500] <= r_data[20499];
                
                r_data[20501] <= r_data[20500];
                
                r_data[20502] <= r_data[20501];
                
                r_data[20503] <= r_data[20502];
                
                r_data[20504] <= r_data[20503];
                
                r_data[20505] <= r_data[20504];
                
                r_data[20506] <= r_data[20505];
                
                r_data[20507] <= r_data[20506];
                
                r_data[20508] <= r_data[20507];
                
                r_data[20509] <= r_data[20508];
                
                r_data[20510] <= r_data[20509];
                
                r_data[20511] <= r_data[20510];
                
                r_data[20512] <= r_data[20511];
                
                r_data[20513] <= r_data[20512];
                
                r_data[20514] <= r_data[20513];
                
                r_data[20515] <= r_data[20514];
                
                r_data[20516] <= r_data[20515];
                
                r_data[20517] <= r_data[20516];
                
                r_data[20518] <= r_data[20517];
                
                r_data[20519] <= r_data[20518];
                
                r_data[20520] <= r_data[20519];
                
                r_data[20521] <= r_data[20520];
                
                r_data[20522] <= r_data[20521];
                
                r_data[20523] <= r_data[20522];
                
                r_data[20524] <= r_data[20523];
                
                r_data[20525] <= r_data[20524];
                
                r_data[20526] <= r_data[20525];
                
                r_data[20527] <= r_data[20526];
                
                r_data[20528] <= r_data[20527];
                
                r_data[20529] <= r_data[20528];
                
                r_data[20530] <= r_data[20529];
                
                r_data[20531] <= r_data[20530];
                
                r_data[20532] <= r_data[20531];
                
                r_data[20533] <= r_data[20532];
                
                r_data[20534] <= r_data[20533];
                
                r_data[20535] <= r_data[20534];
                
                r_data[20536] <= r_data[20535];
                
                r_data[20537] <= r_data[20536];
                
                r_data[20538] <= r_data[20537];
                
                r_data[20539] <= r_data[20538];
                
                r_data[20540] <= r_data[20539];
                
                r_data[20541] <= r_data[20540];
                
                r_data[20542] <= r_data[20541];
                
                r_data[20543] <= r_data[20542];
                
                r_data[20544] <= r_data[20543];
                
                r_data[20545] <= r_data[20544];
                
                r_data[20546] <= r_data[20545];
                
                r_data[20547] <= r_data[20546];
                
                r_data[20548] <= r_data[20547];
                
                r_data[20549] <= r_data[20548];
                
                r_data[20550] <= r_data[20549];
                
                r_data[20551] <= r_data[20550];
                
                r_data[20552] <= r_data[20551];
                
                r_data[20553] <= r_data[20552];
                
                r_data[20554] <= r_data[20553];
                
                r_data[20555] <= r_data[20554];
                
                r_data[20556] <= r_data[20555];
                
                r_data[20557] <= r_data[20556];
                
                r_data[20558] <= r_data[20557];
                
                r_data[20559] <= r_data[20558];
                
                r_data[20560] <= r_data[20559];
                
                r_data[20561] <= r_data[20560];
                
                r_data[20562] <= r_data[20561];
                
                r_data[20563] <= r_data[20562];
                
                r_data[20564] <= r_data[20563];
                
                r_data[20565] <= r_data[20564];
                
                r_data[20566] <= r_data[20565];
                
                r_data[20567] <= r_data[20566];
                
                r_data[20568] <= r_data[20567];
                
                r_data[20569] <= r_data[20568];
                
                r_data[20570] <= r_data[20569];
                
                r_data[20571] <= r_data[20570];
                
                r_data[20572] <= r_data[20571];
                
                r_data[20573] <= r_data[20572];
                
                r_data[20574] <= r_data[20573];
                
                r_data[20575] <= r_data[20574];
                
                r_data[20576] <= r_data[20575];
                
                r_data[20577] <= r_data[20576];
                
                r_data[20578] <= r_data[20577];
                
                r_data[20579] <= r_data[20578];
                
                r_data[20580] <= r_data[20579];
                
                r_data[20581] <= r_data[20580];
                
                r_data[20582] <= r_data[20581];
                
                r_data[20583] <= r_data[20582];
                
                r_data[20584] <= r_data[20583];
                
                r_data[20585] <= r_data[20584];
                
                r_data[20586] <= r_data[20585];
                
                r_data[20587] <= r_data[20586];
                
                r_data[20588] <= r_data[20587];
                
                r_data[20589] <= r_data[20588];
                
                r_data[20590] <= r_data[20589];
                
                r_data[20591] <= r_data[20590];
                
                r_data[20592] <= r_data[20591];
                
                r_data[20593] <= r_data[20592];
                
                r_data[20594] <= r_data[20593];
                
                r_data[20595] <= r_data[20594];
                
                r_data[20596] <= r_data[20595];
                
                r_data[20597] <= r_data[20596];
                
                r_data[20598] <= r_data[20597];
                
                r_data[20599] <= r_data[20598];
                
                r_data[20600] <= r_data[20599];
                
                r_data[20601] <= r_data[20600];
                
                r_data[20602] <= r_data[20601];
                
                r_data[20603] <= r_data[20602];
                
                r_data[20604] <= r_data[20603];
                
                r_data[20605] <= r_data[20604];
                
                r_data[20606] <= r_data[20605];
                
                r_data[20607] <= r_data[20606];
                
                r_data[20608] <= r_data[20607];
                
                r_data[20609] <= r_data[20608];
                
                r_data[20610] <= r_data[20609];
                
                r_data[20611] <= r_data[20610];
                
                r_data[20612] <= r_data[20611];
                
                r_data[20613] <= r_data[20612];
                
                r_data[20614] <= r_data[20613];
                
                r_data[20615] <= r_data[20614];
                
                r_data[20616] <= r_data[20615];
                
                r_data[20617] <= r_data[20616];
                
                r_data[20618] <= r_data[20617];
                
                r_data[20619] <= r_data[20618];
                
                r_data[20620] <= r_data[20619];
                
                r_data[20621] <= r_data[20620];
                
                r_data[20622] <= r_data[20621];
                
                r_data[20623] <= r_data[20622];
                
                r_data[20624] <= r_data[20623];
                
                r_data[20625] <= r_data[20624];
                
                r_data[20626] <= r_data[20625];
                
                r_data[20627] <= r_data[20626];
                
                r_data[20628] <= r_data[20627];
                
                r_data[20629] <= r_data[20628];
                
                r_data[20630] <= r_data[20629];
                
                r_data[20631] <= r_data[20630];
                
                r_data[20632] <= r_data[20631];
                
                r_data[20633] <= r_data[20632];
                
                r_data[20634] <= r_data[20633];
                
                r_data[20635] <= r_data[20634];
                
                r_data[20636] <= r_data[20635];
                
                r_data[20637] <= r_data[20636];
                
                r_data[20638] <= r_data[20637];
                
                r_data[20639] <= r_data[20638];
                
                r_data[20640] <= r_data[20639];
                
                r_data[20641] <= r_data[20640];
                
                r_data[20642] <= r_data[20641];
                
                r_data[20643] <= r_data[20642];
                
                r_data[20644] <= r_data[20643];
                
                r_data[20645] <= r_data[20644];
                
                r_data[20646] <= r_data[20645];
                
                r_data[20647] <= r_data[20646];
                
                r_data[20648] <= r_data[20647];
                
                r_data[20649] <= r_data[20648];
                
                r_data[20650] <= r_data[20649];
                
                r_data[20651] <= r_data[20650];
                
                r_data[20652] <= r_data[20651];
                
                r_data[20653] <= r_data[20652];
                
                r_data[20654] <= r_data[20653];
                
                r_data[20655] <= r_data[20654];
                
                r_data[20656] <= r_data[20655];
                
                r_data[20657] <= r_data[20656];
                
                r_data[20658] <= r_data[20657];
                
                r_data[20659] <= r_data[20658];
                
                r_data[20660] <= r_data[20659];
                
                r_data[20661] <= r_data[20660];
                
                r_data[20662] <= r_data[20661];
                
                r_data[20663] <= r_data[20662];
                
                r_data[20664] <= r_data[20663];
                
                r_data[20665] <= r_data[20664];
                
                r_data[20666] <= r_data[20665];
                
                r_data[20667] <= r_data[20666];
                
                r_data[20668] <= r_data[20667];
                
                r_data[20669] <= r_data[20668];
                
                r_data[20670] <= r_data[20669];
                
                r_data[20671] <= r_data[20670];
                
                r_data[20672] <= r_data[20671];
                
                r_data[20673] <= r_data[20672];
                
                r_data[20674] <= r_data[20673];
                
                r_data[20675] <= r_data[20674];
                
                r_data[20676] <= r_data[20675];
                
                r_data[20677] <= r_data[20676];
                
                r_data[20678] <= r_data[20677];
                
                r_data[20679] <= r_data[20678];
                
                r_data[20680] <= r_data[20679];
                
                r_data[20681] <= r_data[20680];
                
                r_data[20682] <= r_data[20681];
                
                r_data[20683] <= r_data[20682];
                
                r_data[20684] <= r_data[20683];
                
                r_data[20685] <= r_data[20684];
                
                r_data[20686] <= r_data[20685];
                
                r_data[20687] <= r_data[20686];
                
                r_data[20688] <= r_data[20687];
                
                r_data[20689] <= r_data[20688];
                
                r_data[20690] <= r_data[20689];
                
                r_data[20691] <= r_data[20690];
                
                r_data[20692] <= r_data[20691];
                
                r_data[20693] <= r_data[20692];
                
                r_data[20694] <= r_data[20693];
                
                r_data[20695] <= r_data[20694];
                
                r_data[20696] <= r_data[20695];
                
                r_data[20697] <= r_data[20696];
                
                r_data[20698] <= r_data[20697];
                
                r_data[20699] <= r_data[20698];
                
                r_data[20700] <= r_data[20699];
                
                r_data[20701] <= r_data[20700];
                
                r_data[20702] <= r_data[20701];
                
                r_data[20703] <= r_data[20702];
                
                r_data[20704] <= r_data[20703];
                
                r_data[20705] <= r_data[20704];
                
                r_data[20706] <= r_data[20705];
                
                r_data[20707] <= r_data[20706];
                
                r_data[20708] <= r_data[20707];
                
                r_data[20709] <= r_data[20708];
                
                r_data[20710] <= r_data[20709];
                
                r_data[20711] <= r_data[20710];
                
                r_data[20712] <= r_data[20711];
                
                r_data[20713] <= r_data[20712];
                
                r_data[20714] <= r_data[20713];
                
                r_data[20715] <= r_data[20714];
                
                r_data[20716] <= r_data[20715];
                
                r_data[20717] <= r_data[20716];
                
                r_data[20718] <= r_data[20717];
                
                r_data[20719] <= r_data[20718];
                
                r_data[20720] <= r_data[20719];
                
                r_data[20721] <= r_data[20720];
                
                r_data[20722] <= r_data[20721];
                
                r_data[20723] <= r_data[20722];
                
                r_data[20724] <= r_data[20723];
                
                r_data[20725] <= r_data[20724];
                
                r_data[20726] <= r_data[20725];
                
                r_data[20727] <= r_data[20726];
                
                r_data[20728] <= r_data[20727];
                
                r_data[20729] <= r_data[20728];
                
                r_data[20730] <= r_data[20729];
                
                r_data[20731] <= r_data[20730];
                
                r_data[20732] <= r_data[20731];
                
                r_data[20733] <= r_data[20732];
                
                r_data[20734] <= r_data[20733];
                
                r_data[20735] <= r_data[20734];
                
                r_data[20736] <= r_data[20735];
                
                r_data[20737] <= r_data[20736];
                
                r_data[20738] <= r_data[20737];
                
                r_data[20739] <= r_data[20738];
                
                r_data[20740] <= r_data[20739];
                
                r_data[20741] <= r_data[20740];
                
                r_data[20742] <= r_data[20741];
                
                r_data[20743] <= r_data[20742];
                
                r_data[20744] <= r_data[20743];
                
                r_data[20745] <= r_data[20744];
                
                r_data[20746] <= r_data[20745];
                
                r_data[20747] <= r_data[20746];
                
                r_data[20748] <= r_data[20747];
                
                r_data[20749] <= r_data[20748];
                
                r_data[20750] <= r_data[20749];
                
                r_data[20751] <= r_data[20750];
                
                r_data[20752] <= r_data[20751];
                
                r_data[20753] <= r_data[20752];
                
                r_data[20754] <= r_data[20753];
                
                r_data[20755] <= r_data[20754];
                
                r_data[20756] <= r_data[20755];
                
                r_data[20757] <= r_data[20756];
                
                r_data[20758] <= r_data[20757];
                
                r_data[20759] <= r_data[20758];
                
                r_data[20760] <= r_data[20759];
                
                r_data[20761] <= r_data[20760];
                
                r_data[20762] <= r_data[20761];
                
                r_data[20763] <= r_data[20762];
                
                r_data[20764] <= r_data[20763];
                
                r_data[20765] <= r_data[20764];
                
                r_data[20766] <= r_data[20765];
                
                r_data[20767] <= r_data[20766];
                
                r_data[20768] <= r_data[20767];
                
                r_data[20769] <= r_data[20768];
                
                r_data[20770] <= r_data[20769];
                
                r_data[20771] <= r_data[20770];
                
                r_data[20772] <= r_data[20771];
                
                r_data[20773] <= r_data[20772];
                
                r_data[20774] <= r_data[20773];
                
                r_data[20775] <= r_data[20774];
                
                r_data[20776] <= r_data[20775];
                
                r_data[20777] <= r_data[20776];
                
                r_data[20778] <= r_data[20777];
                
                r_data[20779] <= r_data[20778];
                
                r_data[20780] <= r_data[20779];
                
                r_data[20781] <= r_data[20780];
                
                r_data[20782] <= r_data[20781];
                
                r_data[20783] <= r_data[20782];
                
                r_data[20784] <= r_data[20783];
                
                r_data[20785] <= r_data[20784];
                
                r_data[20786] <= r_data[20785];
                
                r_data[20787] <= r_data[20786];
                
                r_data[20788] <= r_data[20787];
                
                r_data[20789] <= r_data[20788];
                
                r_data[20790] <= r_data[20789];
                
                r_data[20791] <= r_data[20790];
                
                r_data[20792] <= r_data[20791];
                
                r_data[20793] <= r_data[20792];
                
                r_data[20794] <= r_data[20793];
                
                r_data[20795] <= r_data[20794];
                
                r_data[20796] <= r_data[20795];
                
                r_data[20797] <= r_data[20796];
                
                r_data[20798] <= r_data[20797];
                
                r_data[20799] <= r_data[20798];
                
                r_data[20800] <= r_data[20799];
                
                r_data[20801] <= r_data[20800];
                
                r_data[20802] <= r_data[20801];
                
                r_data[20803] <= r_data[20802];
                
                r_data[20804] <= r_data[20803];
                
                r_data[20805] <= r_data[20804];
                
                r_data[20806] <= r_data[20805];
                
                r_data[20807] <= r_data[20806];
                
                r_data[20808] <= r_data[20807];
                
                r_data[20809] <= r_data[20808];
                
                r_data[20810] <= r_data[20809];
                
                r_data[20811] <= r_data[20810];
                
                r_data[20812] <= r_data[20811];
                
                r_data[20813] <= r_data[20812];
                
                r_data[20814] <= r_data[20813];
                
                r_data[20815] <= r_data[20814];
                
                r_data[20816] <= r_data[20815];
                
                r_data[20817] <= r_data[20816];
                
                r_data[20818] <= r_data[20817];
                
                r_data[20819] <= r_data[20818];
                
                r_data[20820] <= r_data[20819];
                
                r_data[20821] <= r_data[20820];
                
                r_data[20822] <= r_data[20821];
                
                r_data[20823] <= r_data[20822];
                
                r_data[20824] <= r_data[20823];
                
                r_data[20825] <= r_data[20824];
                
                r_data[20826] <= r_data[20825];
                
                r_data[20827] <= r_data[20826];
                
                r_data[20828] <= r_data[20827];
                
                r_data[20829] <= r_data[20828];
                
                r_data[20830] <= r_data[20829];
                
                r_data[20831] <= r_data[20830];
                
                r_data[20832] <= r_data[20831];
                
                r_data[20833] <= r_data[20832];
                
                r_data[20834] <= r_data[20833];
                
                r_data[20835] <= r_data[20834];
                
                r_data[20836] <= r_data[20835];
                
                r_data[20837] <= r_data[20836];
                
                r_data[20838] <= r_data[20837];
                
                r_data[20839] <= r_data[20838];
                
                r_data[20840] <= r_data[20839];
                
                r_data[20841] <= r_data[20840];
                
                r_data[20842] <= r_data[20841];
                
                r_data[20843] <= r_data[20842];
                
                r_data[20844] <= r_data[20843];
                
                r_data[20845] <= r_data[20844];
                
                r_data[20846] <= r_data[20845];
                
                r_data[20847] <= r_data[20846];
                
                r_data[20848] <= r_data[20847];
                
                r_data[20849] <= r_data[20848];
                
                r_data[20850] <= r_data[20849];
                
                r_data[20851] <= r_data[20850];
                
                r_data[20852] <= r_data[20851];
                
                r_data[20853] <= r_data[20852];
                
                r_data[20854] <= r_data[20853];
                
                r_data[20855] <= r_data[20854];
                
                r_data[20856] <= r_data[20855];
                
                r_data[20857] <= r_data[20856];
                
                r_data[20858] <= r_data[20857];
                
                r_data[20859] <= r_data[20858];
                
                r_data[20860] <= r_data[20859];
                
                r_data[20861] <= r_data[20860];
                
                r_data[20862] <= r_data[20861];
                
                r_data[20863] <= r_data[20862];
                
                r_data[20864] <= r_data[20863];
                
                r_data[20865] <= r_data[20864];
                
                r_data[20866] <= r_data[20865];
                
                r_data[20867] <= r_data[20866];
                
                r_data[20868] <= r_data[20867];
                
                r_data[20869] <= r_data[20868];
                
                r_data[20870] <= r_data[20869];
                
                r_data[20871] <= r_data[20870];
                
                r_data[20872] <= r_data[20871];
                
                r_data[20873] <= r_data[20872];
                
                r_data[20874] <= r_data[20873];
                
                r_data[20875] <= r_data[20874];
                
                r_data[20876] <= r_data[20875];
                
                r_data[20877] <= r_data[20876];
                
                r_data[20878] <= r_data[20877];
                
                r_data[20879] <= r_data[20878];
                
                r_data[20880] <= r_data[20879];
                
                r_data[20881] <= r_data[20880];
                
                r_data[20882] <= r_data[20881];
                
                r_data[20883] <= r_data[20882];
                
                r_data[20884] <= r_data[20883];
                
                r_data[20885] <= r_data[20884];
                
                r_data[20886] <= r_data[20885];
                
                r_data[20887] <= r_data[20886];
                
                r_data[20888] <= r_data[20887];
                
                r_data[20889] <= r_data[20888];
                
                r_data[20890] <= r_data[20889];
                
                r_data[20891] <= r_data[20890];
                
                r_data[20892] <= r_data[20891];
                
                r_data[20893] <= r_data[20892];
                
                r_data[20894] <= r_data[20893];
                
                r_data[20895] <= r_data[20894];
                
                r_data[20896] <= r_data[20895];
                
                r_data[20897] <= r_data[20896];
                
                r_data[20898] <= r_data[20897];
                
                r_data[20899] <= r_data[20898];
                
                r_data[20900] <= r_data[20899];
                
                r_data[20901] <= r_data[20900];
                
                r_data[20902] <= r_data[20901];
                
                r_data[20903] <= r_data[20902];
                
                r_data[20904] <= r_data[20903];
                
                r_data[20905] <= r_data[20904];
                
                r_data[20906] <= r_data[20905];
                
                r_data[20907] <= r_data[20906];
                
                r_data[20908] <= r_data[20907];
                
                r_data[20909] <= r_data[20908];
                
                r_data[20910] <= r_data[20909];
                
                r_data[20911] <= r_data[20910];
                
                r_data[20912] <= r_data[20911];
                
                r_data[20913] <= r_data[20912];
                
                r_data[20914] <= r_data[20913];
                
                r_data[20915] <= r_data[20914];
                
                r_data[20916] <= r_data[20915];
                
                r_data[20917] <= r_data[20916];
                
                r_data[20918] <= r_data[20917];
                
                r_data[20919] <= r_data[20918];
                
                r_data[20920] <= r_data[20919];
                
                r_data[20921] <= r_data[20920];
                
                r_data[20922] <= r_data[20921];
                
                r_data[20923] <= r_data[20922];
                
                r_data[20924] <= r_data[20923];
                
                r_data[20925] <= r_data[20924];
                
                r_data[20926] <= r_data[20925];
                
                r_data[20927] <= r_data[20926];
                
                r_data[20928] <= r_data[20927];
                
                r_data[20929] <= r_data[20928];
                
                r_data[20930] <= r_data[20929];
                
                r_data[20931] <= r_data[20930];
                
                r_data[20932] <= r_data[20931];
                
                r_data[20933] <= r_data[20932];
                
                r_data[20934] <= r_data[20933];
                
                r_data[20935] <= r_data[20934];
                
                r_data[20936] <= r_data[20935];
                
                r_data[20937] <= r_data[20936];
                
                r_data[20938] <= r_data[20937];
                
                r_data[20939] <= r_data[20938];
                
                r_data[20940] <= r_data[20939];
                
                r_data[20941] <= r_data[20940];
                
                r_data[20942] <= r_data[20941];
                
                r_data[20943] <= r_data[20942];
                
                r_data[20944] <= r_data[20943];
                
                r_data[20945] <= r_data[20944];
                
                r_data[20946] <= r_data[20945];
                
                r_data[20947] <= r_data[20946];
                
                r_data[20948] <= r_data[20947];
                
                r_data[20949] <= r_data[20948];
                
                r_data[20950] <= r_data[20949];
                
                r_data[20951] <= r_data[20950];
                
                r_data[20952] <= r_data[20951];
                
                r_data[20953] <= r_data[20952];
                
                r_data[20954] <= r_data[20953];
                
                r_data[20955] <= r_data[20954];
                
                r_data[20956] <= r_data[20955];
                
                r_data[20957] <= r_data[20956];
                
                r_data[20958] <= r_data[20957];
                
                r_data[20959] <= r_data[20958];
                
                r_data[20960] <= r_data[20959];
                
                r_data[20961] <= r_data[20960];
                
                r_data[20962] <= r_data[20961];
                
                r_data[20963] <= r_data[20962];
                
                r_data[20964] <= r_data[20963];
                
                r_data[20965] <= r_data[20964];
                
                r_data[20966] <= r_data[20965];
                
                r_data[20967] <= r_data[20966];
                
                r_data[20968] <= r_data[20967];
                
                r_data[20969] <= r_data[20968];
                
                r_data[20970] <= r_data[20969];
                
                r_data[20971] <= r_data[20970];
                
                r_data[20972] <= r_data[20971];
                
                r_data[20973] <= r_data[20972];
                
                r_data[20974] <= r_data[20973];
                
                r_data[20975] <= r_data[20974];
                
                r_data[20976] <= r_data[20975];
                
                r_data[20977] <= r_data[20976];
                
                r_data[20978] <= r_data[20977];
                
                r_data[20979] <= r_data[20978];
                
                r_data[20980] <= r_data[20979];
                
                r_data[20981] <= r_data[20980];
                
                r_data[20982] <= r_data[20981];
                
                r_data[20983] <= r_data[20982];
                
                r_data[20984] <= r_data[20983];
                
                r_data[20985] <= r_data[20984];
                
                r_data[20986] <= r_data[20985];
                
                r_data[20987] <= r_data[20986];
                
                r_data[20988] <= r_data[20987];
                
                r_data[20989] <= r_data[20988];
                
                r_data[20990] <= r_data[20989];
                
                r_data[20991] <= r_data[20990];
                
                r_data[20992] <= r_data[20991];
                
                r_data[20993] <= r_data[20992];
                
                r_data[20994] <= r_data[20993];
                
                r_data[20995] <= r_data[20994];
                
                r_data[20996] <= r_data[20995];
                
                r_data[20997] <= r_data[20996];
                
                r_data[20998] <= r_data[20997];
                
                r_data[20999] <= r_data[20998];
                
                r_data[21000] <= r_data[20999];
                
                r_data[21001] <= r_data[21000];
                
                r_data[21002] <= r_data[21001];
                
                r_data[21003] <= r_data[21002];
                
                r_data[21004] <= r_data[21003];
                
                r_data[21005] <= r_data[21004];
                
                r_data[21006] <= r_data[21005];
                
                r_data[21007] <= r_data[21006];
                
                r_data[21008] <= r_data[21007];
                
                r_data[21009] <= r_data[21008];
                
                r_data[21010] <= r_data[21009];
                
                r_data[21011] <= r_data[21010];
                
                r_data[21012] <= r_data[21011];
                
                r_data[21013] <= r_data[21012];
                
                r_data[21014] <= r_data[21013];
                
                r_data[21015] <= r_data[21014];
                
                r_data[21016] <= r_data[21015];
                
                r_data[21017] <= r_data[21016];
                
                r_data[21018] <= r_data[21017];
                
                r_data[21019] <= r_data[21018];
                
                r_data[21020] <= r_data[21019];
                
                r_data[21021] <= r_data[21020];
                
                r_data[21022] <= r_data[21021];
                
                r_data[21023] <= r_data[21022];
                
                r_data[21024] <= r_data[21023];
                
                r_data[21025] <= r_data[21024];
                
                r_data[21026] <= r_data[21025];
                
                r_data[21027] <= r_data[21026];
                
                r_data[21028] <= r_data[21027];
                
                r_data[21029] <= r_data[21028];
                
                r_data[21030] <= r_data[21029];
                
                r_data[21031] <= r_data[21030];
                
                r_data[21032] <= r_data[21031];
                
                r_data[21033] <= r_data[21032];
                
                r_data[21034] <= r_data[21033];
                
                r_data[21035] <= r_data[21034];
                
                r_data[21036] <= r_data[21035];
                
                r_data[21037] <= r_data[21036];
                
                r_data[21038] <= r_data[21037];
                
                r_data[21039] <= r_data[21038];
                
                r_data[21040] <= r_data[21039];
                
                r_data[21041] <= r_data[21040];
                
                r_data[21042] <= r_data[21041];
                
                r_data[21043] <= r_data[21042];
                
                r_data[21044] <= r_data[21043];
                
                r_data[21045] <= r_data[21044];
                
                r_data[21046] <= r_data[21045];
                
                r_data[21047] <= r_data[21046];
                
                r_data[21048] <= r_data[21047];
                
                r_data[21049] <= r_data[21048];
                
                r_data[21050] <= r_data[21049];
                
                r_data[21051] <= r_data[21050];
                
                r_data[21052] <= r_data[21051];
                
                r_data[21053] <= r_data[21052];
                
                r_data[21054] <= r_data[21053];
                
                r_data[21055] <= r_data[21054];
                
                r_data[21056] <= r_data[21055];
                
                r_data[21057] <= r_data[21056];
                
                r_data[21058] <= r_data[21057];
                
                r_data[21059] <= r_data[21058];
                
                r_data[21060] <= r_data[21059];
                
                r_data[21061] <= r_data[21060];
                
                r_data[21062] <= r_data[21061];
                
                r_data[21063] <= r_data[21062];
                
                r_data[21064] <= r_data[21063];
                
                r_data[21065] <= r_data[21064];
                
                r_data[21066] <= r_data[21065];
                
                r_data[21067] <= r_data[21066];
                
                r_data[21068] <= r_data[21067];
                
                r_data[21069] <= r_data[21068];
                
                r_data[21070] <= r_data[21069];
                
                r_data[21071] <= r_data[21070];
                
                r_data[21072] <= r_data[21071];
                
                r_data[21073] <= r_data[21072];
                
                r_data[21074] <= r_data[21073];
                
                r_data[21075] <= r_data[21074];
                
                r_data[21076] <= r_data[21075];
                
                r_data[21077] <= r_data[21076];
                
                r_data[21078] <= r_data[21077];
                
                r_data[21079] <= r_data[21078];
                
                r_data[21080] <= r_data[21079];
                
                r_data[21081] <= r_data[21080];
                
                r_data[21082] <= r_data[21081];
                
                r_data[21083] <= r_data[21082];
                
                r_data[21084] <= r_data[21083];
                
                r_data[21085] <= r_data[21084];
                
                r_data[21086] <= r_data[21085];
                
                r_data[21087] <= r_data[21086];
                
                r_data[21088] <= r_data[21087];
                
                r_data[21089] <= r_data[21088];
                
                r_data[21090] <= r_data[21089];
                
                r_data[21091] <= r_data[21090];
                
                r_data[21092] <= r_data[21091];
                
                r_data[21093] <= r_data[21092];
                
                r_data[21094] <= r_data[21093];
                
                r_data[21095] <= r_data[21094];
                
                r_data[21096] <= r_data[21095];
                
                r_data[21097] <= r_data[21096];
                
                r_data[21098] <= r_data[21097];
                
                r_data[21099] <= r_data[21098];
                
                r_data[21100] <= r_data[21099];
                
                r_data[21101] <= r_data[21100];
                
                r_data[21102] <= r_data[21101];
                
                r_data[21103] <= r_data[21102];
                
                r_data[21104] <= r_data[21103];
                
                r_data[21105] <= r_data[21104];
                
                r_data[21106] <= r_data[21105];
                
                r_data[21107] <= r_data[21106];
                
                r_data[21108] <= r_data[21107];
                
                r_data[21109] <= r_data[21108];
                
                r_data[21110] <= r_data[21109];
                
                r_data[21111] <= r_data[21110];
                
                r_data[21112] <= r_data[21111];
                
                r_data[21113] <= r_data[21112];
                
                r_data[21114] <= r_data[21113];
                
                r_data[21115] <= r_data[21114];
                
                r_data[21116] <= r_data[21115];
                
                r_data[21117] <= r_data[21116];
                
                r_data[21118] <= r_data[21117];
                
                r_data[21119] <= r_data[21118];
                
                r_data[21120] <= r_data[21119];
                
                r_data[21121] <= r_data[21120];
                
                r_data[21122] <= r_data[21121];
                
                r_data[21123] <= r_data[21122];
                
                r_data[21124] <= r_data[21123];
                
                r_data[21125] <= r_data[21124];
                
                r_data[21126] <= r_data[21125];
                
                r_data[21127] <= r_data[21126];
                
                r_data[21128] <= r_data[21127];
                
                r_data[21129] <= r_data[21128];
                
                r_data[21130] <= r_data[21129];
                
                r_data[21131] <= r_data[21130];
                
                r_data[21132] <= r_data[21131];
                
                r_data[21133] <= r_data[21132];
                
                r_data[21134] <= r_data[21133];
                
                r_data[21135] <= r_data[21134];
                
                r_data[21136] <= r_data[21135];
                
                r_data[21137] <= r_data[21136];
                
                r_data[21138] <= r_data[21137];
                
                r_data[21139] <= r_data[21138];
                
                r_data[21140] <= r_data[21139];
                
                r_data[21141] <= r_data[21140];
                
                r_data[21142] <= r_data[21141];
                
                r_data[21143] <= r_data[21142];
                
                r_data[21144] <= r_data[21143];
                
                r_data[21145] <= r_data[21144];
                
                r_data[21146] <= r_data[21145];
                
                r_data[21147] <= r_data[21146];
                
                r_data[21148] <= r_data[21147];
                
                r_data[21149] <= r_data[21148];
                
                r_data[21150] <= r_data[21149];
                
                r_data[21151] <= r_data[21150];
                
                r_data[21152] <= r_data[21151];
                
                r_data[21153] <= r_data[21152];
                
                r_data[21154] <= r_data[21153];
                
                r_data[21155] <= r_data[21154];
                
                r_data[21156] <= r_data[21155];
                
                r_data[21157] <= r_data[21156];
                
                r_data[21158] <= r_data[21157];
                
                r_data[21159] <= r_data[21158];
                
                r_data[21160] <= r_data[21159];
                
                r_data[21161] <= r_data[21160];
                
                r_data[21162] <= r_data[21161];
                
                r_data[21163] <= r_data[21162];
                
                r_data[21164] <= r_data[21163];
                
                r_data[21165] <= r_data[21164];
                
                r_data[21166] <= r_data[21165];
                
                r_data[21167] <= r_data[21166];
                
                r_data[21168] <= r_data[21167];
                
                r_data[21169] <= r_data[21168];
                
                r_data[21170] <= r_data[21169];
                
                r_data[21171] <= r_data[21170];
                
                r_data[21172] <= r_data[21171];
                
                r_data[21173] <= r_data[21172];
                
                r_data[21174] <= r_data[21173];
                
                r_data[21175] <= r_data[21174];
                
                r_data[21176] <= r_data[21175];
                
                r_data[21177] <= r_data[21176];
                
                r_data[21178] <= r_data[21177];
                
                r_data[21179] <= r_data[21178];
                
                r_data[21180] <= r_data[21179];
                
                r_data[21181] <= r_data[21180];
                
                r_data[21182] <= r_data[21181];
                
                r_data[21183] <= r_data[21182];
                
                r_data[21184] <= r_data[21183];
                
                r_data[21185] <= r_data[21184];
                
                r_data[21186] <= r_data[21185];
                
                r_data[21187] <= r_data[21186];
                
                r_data[21188] <= r_data[21187];
                
                r_data[21189] <= r_data[21188];
                
                r_data[21190] <= r_data[21189];
                
                r_data[21191] <= r_data[21190];
                
                r_data[21192] <= r_data[21191];
                
                r_data[21193] <= r_data[21192];
                
                r_data[21194] <= r_data[21193];
                
                r_data[21195] <= r_data[21194];
                
                r_data[21196] <= r_data[21195];
                
                r_data[21197] <= r_data[21196];
                
                r_data[21198] <= r_data[21197];
                
                r_data[21199] <= r_data[21198];
                
                r_data[21200] <= r_data[21199];
                
                r_data[21201] <= r_data[21200];
                
                r_data[21202] <= r_data[21201];
                
                r_data[21203] <= r_data[21202];
                
                r_data[21204] <= r_data[21203];
                
                r_data[21205] <= r_data[21204];
                
                r_data[21206] <= r_data[21205];
                
                r_data[21207] <= r_data[21206];
                
                r_data[21208] <= r_data[21207];
                
                r_data[21209] <= r_data[21208];
                
                r_data[21210] <= r_data[21209];
                
                r_data[21211] <= r_data[21210];
                
                r_data[21212] <= r_data[21211];
                
                r_data[21213] <= r_data[21212];
                
                r_data[21214] <= r_data[21213];
                
                r_data[21215] <= r_data[21214];
                
                r_data[21216] <= r_data[21215];
                
                r_data[21217] <= r_data[21216];
                
                r_data[21218] <= r_data[21217];
                
                r_data[21219] <= r_data[21218];
                
                r_data[21220] <= r_data[21219];
                
                r_data[21221] <= r_data[21220];
                
                r_data[21222] <= r_data[21221];
                
                r_data[21223] <= r_data[21222];
                
                r_data[21224] <= r_data[21223];
                
                r_data[21225] <= r_data[21224];
                
                r_data[21226] <= r_data[21225];
                
                r_data[21227] <= r_data[21226];
                
                r_data[21228] <= r_data[21227];
                
                r_data[21229] <= r_data[21228];
                
                r_data[21230] <= r_data[21229];
                
                r_data[21231] <= r_data[21230];
                
                r_data[21232] <= r_data[21231];
                
                r_data[21233] <= r_data[21232];
                
                r_data[21234] <= r_data[21233];
                
                r_data[21235] <= r_data[21234];
                
                r_data[21236] <= r_data[21235];
                
                r_data[21237] <= r_data[21236];
                
                r_data[21238] <= r_data[21237];
                
                r_data[21239] <= r_data[21238];
                
                r_data[21240] <= r_data[21239];
                
                r_data[21241] <= r_data[21240];
                
                r_data[21242] <= r_data[21241];
                
                r_data[21243] <= r_data[21242];
                
                r_data[21244] <= r_data[21243];
                
                r_data[21245] <= r_data[21244];
                
                r_data[21246] <= r_data[21245];
                
                r_data[21247] <= r_data[21246];
                
                r_data[21248] <= r_data[21247];
                
                r_data[21249] <= r_data[21248];
                
                r_data[21250] <= r_data[21249];
                
                r_data[21251] <= r_data[21250];
                
                r_data[21252] <= r_data[21251];
                
                r_data[21253] <= r_data[21252];
                
                r_data[21254] <= r_data[21253];
                
                r_data[21255] <= r_data[21254];
                
                r_data[21256] <= r_data[21255];
                
                r_data[21257] <= r_data[21256];
                
                r_data[21258] <= r_data[21257];
                
                r_data[21259] <= r_data[21258];
                
                r_data[21260] <= r_data[21259];
                
                r_data[21261] <= r_data[21260];
                
                r_data[21262] <= r_data[21261];
                
                r_data[21263] <= r_data[21262];
                
                r_data[21264] <= r_data[21263];
                
                r_data[21265] <= r_data[21264];
                
                r_data[21266] <= r_data[21265];
                
                r_data[21267] <= r_data[21266];
                
                r_data[21268] <= r_data[21267];
                
                r_data[21269] <= r_data[21268];
                
                r_data[21270] <= r_data[21269];
                
                r_data[21271] <= r_data[21270];
                
                r_data[21272] <= r_data[21271];
                
                r_data[21273] <= r_data[21272];
                
                r_data[21274] <= r_data[21273];
                
                r_data[21275] <= r_data[21274];
                
                r_data[21276] <= r_data[21275];
                
                r_data[21277] <= r_data[21276];
                
                r_data[21278] <= r_data[21277];
                
                r_data[21279] <= r_data[21278];
                
                r_data[21280] <= r_data[21279];
                
                r_data[21281] <= r_data[21280];
                
                r_data[21282] <= r_data[21281];
                
                r_data[21283] <= r_data[21282];
                
                r_data[21284] <= r_data[21283];
                
                r_data[21285] <= r_data[21284];
                
                r_data[21286] <= r_data[21285];
                
                r_data[21287] <= r_data[21286];
                
                r_data[21288] <= r_data[21287];
                
                r_data[21289] <= r_data[21288];
                
                r_data[21290] <= r_data[21289];
                
                r_data[21291] <= r_data[21290];
                
                r_data[21292] <= r_data[21291];
                
                r_data[21293] <= r_data[21292];
                
                r_data[21294] <= r_data[21293];
                
                r_data[21295] <= r_data[21294];
                
                r_data[21296] <= r_data[21295];
                
                r_data[21297] <= r_data[21296];
                
                r_data[21298] <= r_data[21297];
                
                r_data[21299] <= r_data[21298];
                
                r_data[21300] <= r_data[21299];
                
                r_data[21301] <= r_data[21300];
                
                r_data[21302] <= r_data[21301];
                
                r_data[21303] <= r_data[21302];
                
                r_data[21304] <= r_data[21303];
                
                r_data[21305] <= r_data[21304];
                
                r_data[21306] <= r_data[21305];
                
                r_data[21307] <= r_data[21306];
                
                r_data[21308] <= r_data[21307];
                
                r_data[21309] <= r_data[21308];
                
                r_data[21310] <= r_data[21309];
                
                r_data[21311] <= r_data[21310];
                
                r_data[21312] <= r_data[21311];
                
                r_data[21313] <= r_data[21312];
                
                r_data[21314] <= r_data[21313];
                
                r_data[21315] <= r_data[21314];
                
                r_data[21316] <= r_data[21315];
                
                r_data[21317] <= r_data[21316];
                
                r_data[21318] <= r_data[21317];
                
                r_data[21319] <= r_data[21318];
                
                r_data[21320] <= r_data[21319];
                
                r_data[21321] <= r_data[21320];
                
                r_data[21322] <= r_data[21321];
                
                r_data[21323] <= r_data[21322];
                
                r_data[21324] <= r_data[21323];
                
                r_data[21325] <= r_data[21324];
                
                r_data[21326] <= r_data[21325];
                
                r_data[21327] <= r_data[21326];
                
                r_data[21328] <= r_data[21327];
                
                r_data[21329] <= r_data[21328];
                
                r_data[21330] <= r_data[21329];
                
                r_data[21331] <= r_data[21330];
                
                r_data[21332] <= r_data[21331];
                
                r_data[21333] <= r_data[21332];
                
                r_data[21334] <= r_data[21333];
                
                r_data[21335] <= r_data[21334];
                
                r_data[21336] <= r_data[21335];
                
                r_data[21337] <= r_data[21336];
                
                r_data[21338] <= r_data[21337];
                
                r_data[21339] <= r_data[21338];
                
                r_data[21340] <= r_data[21339];
                
                r_data[21341] <= r_data[21340];
                
                r_data[21342] <= r_data[21341];
                
                r_data[21343] <= r_data[21342];
                
                r_data[21344] <= r_data[21343];
                
                r_data[21345] <= r_data[21344];
                
                r_data[21346] <= r_data[21345];
                
                r_data[21347] <= r_data[21346];
                
                r_data[21348] <= r_data[21347];
                
                r_data[21349] <= r_data[21348];
                
                r_data[21350] <= r_data[21349];
                
                r_data[21351] <= r_data[21350];
                
                r_data[21352] <= r_data[21351];
                
                r_data[21353] <= r_data[21352];
                
                r_data[21354] <= r_data[21353];
                
                r_data[21355] <= r_data[21354];
                
                r_data[21356] <= r_data[21355];
                
                r_data[21357] <= r_data[21356];
                
                r_data[21358] <= r_data[21357];
                
                r_data[21359] <= r_data[21358];
                
                r_data[21360] <= r_data[21359];
                
                r_data[21361] <= r_data[21360];
                
                r_data[21362] <= r_data[21361];
                
                r_data[21363] <= r_data[21362];
                
                r_data[21364] <= r_data[21363];
                
                r_data[21365] <= r_data[21364];
                
                r_data[21366] <= r_data[21365];
                
                r_data[21367] <= r_data[21366];
                
                r_data[21368] <= r_data[21367];
                
                r_data[21369] <= r_data[21368];
                
                r_data[21370] <= r_data[21369];
                
                r_data[21371] <= r_data[21370];
                
                r_data[21372] <= r_data[21371];
                
                r_data[21373] <= r_data[21372];
                
                r_data[21374] <= r_data[21373];
                
                r_data[21375] <= r_data[21374];
                
                r_data[21376] <= r_data[21375];
                
                r_data[21377] <= r_data[21376];
                
                r_data[21378] <= r_data[21377];
                
                r_data[21379] <= r_data[21378];
                
                r_data[21380] <= r_data[21379];
                
                r_data[21381] <= r_data[21380];
                
                r_data[21382] <= r_data[21381];
                
                r_data[21383] <= r_data[21382];
                
                r_data[21384] <= r_data[21383];
                
                r_data[21385] <= r_data[21384];
                
                r_data[21386] <= r_data[21385];
                
                r_data[21387] <= r_data[21386];
                
                r_data[21388] <= r_data[21387];
                
                r_data[21389] <= r_data[21388];
                
                r_data[21390] <= r_data[21389];
                
                r_data[21391] <= r_data[21390];
                
                r_data[21392] <= r_data[21391];
                
                r_data[21393] <= r_data[21392];
                
                r_data[21394] <= r_data[21393];
                
                r_data[21395] <= r_data[21394];
                
                r_data[21396] <= r_data[21395];
                
                r_data[21397] <= r_data[21396];
                
                r_data[21398] <= r_data[21397];
                
                r_data[21399] <= r_data[21398];
                
                r_data[21400] <= r_data[21399];
                
                r_data[21401] <= r_data[21400];
                
                r_data[21402] <= r_data[21401];
                
                r_data[21403] <= r_data[21402];
                
                r_data[21404] <= r_data[21403];
                
                r_data[21405] <= r_data[21404];
                
                r_data[21406] <= r_data[21405];
                
                r_data[21407] <= r_data[21406];
                
                r_data[21408] <= r_data[21407];
                
                r_data[21409] <= r_data[21408];
                
                r_data[21410] <= r_data[21409];
                
                r_data[21411] <= r_data[21410];
                
                r_data[21412] <= r_data[21411];
                
                r_data[21413] <= r_data[21412];
                
                r_data[21414] <= r_data[21413];
                
                r_data[21415] <= r_data[21414];
                
                r_data[21416] <= r_data[21415];
                
                r_data[21417] <= r_data[21416];
                
                r_data[21418] <= r_data[21417];
                
                r_data[21419] <= r_data[21418];
                
                r_data[21420] <= r_data[21419];
                
                r_data[21421] <= r_data[21420];
                
                r_data[21422] <= r_data[21421];
                
                r_data[21423] <= r_data[21422];
                
                r_data[21424] <= r_data[21423];
                
                r_data[21425] <= r_data[21424];
                
                r_data[21426] <= r_data[21425];
                
                r_data[21427] <= r_data[21426];
                
                r_data[21428] <= r_data[21427];
                
                r_data[21429] <= r_data[21428];
                
                r_data[21430] <= r_data[21429];
                
                r_data[21431] <= r_data[21430];
                
                r_data[21432] <= r_data[21431];
                
                r_data[21433] <= r_data[21432];
                
                r_data[21434] <= r_data[21433];
                
                r_data[21435] <= r_data[21434];
                
                r_data[21436] <= r_data[21435];
                
                r_data[21437] <= r_data[21436];
                
                r_data[21438] <= r_data[21437];
                
                r_data[21439] <= r_data[21438];
                
                r_data[21440] <= r_data[21439];
                
                r_data[21441] <= r_data[21440];
                
                r_data[21442] <= r_data[21441];
                
                r_data[21443] <= r_data[21442];
                
                r_data[21444] <= r_data[21443];
                
                r_data[21445] <= r_data[21444];
                
                r_data[21446] <= r_data[21445];
                
                r_data[21447] <= r_data[21446];
                
                r_data[21448] <= r_data[21447];
                
                r_data[21449] <= r_data[21448];
                
                r_data[21450] <= r_data[21449];
                
                r_data[21451] <= r_data[21450];
                
                r_data[21452] <= r_data[21451];
                
                r_data[21453] <= r_data[21452];
                
                r_data[21454] <= r_data[21453];
                
                r_data[21455] <= r_data[21454];
                
                r_data[21456] <= r_data[21455];
                
                r_data[21457] <= r_data[21456];
                
                r_data[21458] <= r_data[21457];
                
                r_data[21459] <= r_data[21458];
                
                r_data[21460] <= r_data[21459];
                
                r_data[21461] <= r_data[21460];
                
                r_data[21462] <= r_data[21461];
                
                r_data[21463] <= r_data[21462];
                
                r_data[21464] <= r_data[21463];
                
                r_data[21465] <= r_data[21464];
                
                r_data[21466] <= r_data[21465];
                
                r_data[21467] <= r_data[21466];
                
                r_data[21468] <= r_data[21467];
                
                r_data[21469] <= r_data[21468];
                
                r_data[21470] <= r_data[21469];
                
                r_data[21471] <= r_data[21470];
                
                r_data[21472] <= r_data[21471];
                
                r_data[21473] <= r_data[21472];
                
                r_data[21474] <= r_data[21473];
                
                r_data[21475] <= r_data[21474];
                
                r_data[21476] <= r_data[21475];
                
                r_data[21477] <= r_data[21476];
                
                r_data[21478] <= r_data[21477];
                
                r_data[21479] <= r_data[21478];
                
                r_data[21480] <= r_data[21479];
                
                r_data[21481] <= r_data[21480];
                
                r_data[21482] <= r_data[21481];
                
                r_data[21483] <= r_data[21482];
                
                r_data[21484] <= r_data[21483];
                
                r_data[21485] <= r_data[21484];
                
                r_data[21486] <= r_data[21485];
                
                r_data[21487] <= r_data[21486];
                
                r_data[21488] <= r_data[21487];
                
                r_data[21489] <= r_data[21488];
                
                r_data[21490] <= r_data[21489];
                
                r_data[21491] <= r_data[21490];
                
                r_data[21492] <= r_data[21491];
                
                r_data[21493] <= r_data[21492];
                
                r_data[21494] <= r_data[21493];
                
                r_data[21495] <= r_data[21494];
                
                r_data[21496] <= r_data[21495];
                
                r_data[21497] <= r_data[21496];
                
                r_data[21498] <= r_data[21497];
                
                r_data[21499] <= r_data[21498];
                
                r_data[21500] <= r_data[21499];
                
                r_data[21501] <= r_data[21500];
                
                r_data[21502] <= r_data[21501];
                
                r_data[21503] <= r_data[21502];
                
                r_data[21504] <= r_data[21503];
                
                r_data[21505] <= r_data[21504];
                
                r_data[21506] <= r_data[21505];
                
                r_data[21507] <= r_data[21506];
                
                r_data[21508] <= r_data[21507];
                
                r_data[21509] <= r_data[21508];
                
                r_data[21510] <= r_data[21509];
                
                r_data[21511] <= r_data[21510];
                
                r_data[21512] <= r_data[21511];
                
                r_data[21513] <= r_data[21512];
                
                r_data[21514] <= r_data[21513];
                
                r_data[21515] <= r_data[21514];
                
                r_data[21516] <= r_data[21515];
                
                r_data[21517] <= r_data[21516];
                
                r_data[21518] <= r_data[21517];
                
                r_data[21519] <= r_data[21518];
                
                r_data[21520] <= r_data[21519];
                
                r_data[21521] <= r_data[21520];
                
                r_data[21522] <= r_data[21521];
                
                r_data[21523] <= r_data[21522];
                
                r_data[21524] <= r_data[21523];
                
                r_data[21525] <= r_data[21524];
                
                r_data[21526] <= r_data[21525];
                
                r_data[21527] <= r_data[21526];
                
                r_data[21528] <= r_data[21527];
                
                r_data[21529] <= r_data[21528];
                
                r_data[21530] <= r_data[21529];
                
                r_data[21531] <= r_data[21530];
                
                r_data[21532] <= r_data[21531];
                
                r_data[21533] <= r_data[21532];
                
                r_data[21534] <= r_data[21533];
                
                r_data[21535] <= r_data[21534];
                
                r_data[21536] <= r_data[21535];
                
                r_data[21537] <= r_data[21536];
                
                r_data[21538] <= r_data[21537];
                
                r_data[21539] <= r_data[21538];
                
                r_data[21540] <= r_data[21539];
                
                r_data[21541] <= r_data[21540];
                
                r_data[21542] <= r_data[21541];
                
                r_data[21543] <= r_data[21542];
                
                r_data[21544] <= r_data[21543];
                
                r_data[21545] <= r_data[21544];
                
                r_data[21546] <= r_data[21545];
                
                r_data[21547] <= r_data[21546];
                
                r_data[21548] <= r_data[21547];
                
                r_data[21549] <= r_data[21548];
                
                r_data[21550] <= r_data[21549];
                
                r_data[21551] <= r_data[21550];
                
                r_data[21552] <= r_data[21551];
                
                r_data[21553] <= r_data[21552];
                
                r_data[21554] <= r_data[21553];
                
                r_data[21555] <= r_data[21554];
                
                r_data[21556] <= r_data[21555];
                
                r_data[21557] <= r_data[21556];
                
                r_data[21558] <= r_data[21557];
                
                r_data[21559] <= r_data[21558];
                
                r_data[21560] <= r_data[21559];
                
                r_data[21561] <= r_data[21560];
                
                r_data[21562] <= r_data[21561];
                
                r_data[21563] <= r_data[21562];
                
                r_data[21564] <= r_data[21563];
                
                r_data[21565] <= r_data[21564];
                
                r_data[21566] <= r_data[21565];
                
                r_data[21567] <= r_data[21566];
                
                r_data[21568] <= r_data[21567];
                
                r_data[21569] <= r_data[21568];
                
                r_data[21570] <= r_data[21569];
                
                r_data[21571] <= r_data[21570];
                
                r_data[21572] <= r_data[21571];
                
                r_data[21573] <= r_data[21572];
                
                r_data[21574] <= r_data[21573];
                
                r_data[21575] <= r_data[21574];
                
                r_data[21576] <= r_data[21575];
                
                r_data[21577] <= r_data[21576];
                
                r_data[21578] <= r_data[21577];
                
                r_data[21579] <= r_data[21578];
                
                r_data[21580] <= r_data[21579];
                
                r_data[21581] <= r_data[21580];
                
                r_data[21582] <= r_data[21581];
                
                r_data[21583] <= r_data[21582];
                
                r_data[21584] <= r_data[21583];
                
                r_data[21585] <= r_data[21584];
                
                r_data[21586] <= r_data[21585];
                
                r_data[21587] <= r_data[21586];
                
                r_data[21588] <= r_data[21587];
                
                r_data[21589] <= r_data[21588];
                
                r_data[21590] <= r_data[21589];
                
                r_data[21591] <= r_data[21590];
                
                r_data[21592] <= r_data[21591];
                
                r_data[21593] <= r_data[21592];
                
                r_data[21594] <= r_data[21593];
                
                r_data[21595] <= r_data[21594];
                
                r_data[21596] <= r_data[21595];
                
                r_data[21597] <= r_data[21596];
                
                r_data[21598] <= r_data[21597];
                
                r_data[21599] <= r_data[21598];
                
                r_data[21600] <= r_data[21599];
                
                r_data[21601] <= r_data[21600];
                
                r_data[21602] <= r_data[21601];
                
                r_data[21603] <= r_data[21602];
                
                r_data[21604] <= r_data[21603];
                
                r_data[21605] <= r_data[21604];
                
                r_data[21606] <= r_data[21605];
                
                r_data[21607] <= r_data[21606];
                
                r_data[21608] <= r_data[21607];
                
                r_data[21609] <= r_data[21608];
                
                r_data[21610] <= r_data[21609];
                
                r_data[21611] <= r_data[21610];
                
                r_data[21612] <= r_data[21611];
                
                r_data[21613] <= r_data[21612];
                
                r_data[21614] <= r_data[21613];
                
                r_data[21615] <= r_data[21614];
                
                r_data[21616] <= r_data[21615];
                
                r_data[21617] <= r_data[21616];
                
                r_data[21618] <= r_data[21617];
                
                r_data[21619] <= r_data[21618];
                
                r_data[21620] <= r_data[21619];
                
                r_data[21621] <= r_data[21620];
                
                r_data[21622] <= r_data[21621];
                
                r_data[21623] <= r_data[21622];
                
                r_data[21624] <= r_data[21623];
                
                r_data[21625] <= r_data[21624];
                
                r_data[21626] <= r_data[21625];
                
                r_data[21627] <= r_data[21626];
                
                r_data[21628] <= r_data[21627];
                
                r_data[21629] <= r_data[21628];
                
                r_data[21630] <= r_data[21629];
                
                r_data[21631] <= r_data[21630];
                
                r_data[21632] <= r_data[21631];
                
                r_data[21633] <= r_data[21632];
                
                r_data[21634] <= r_data[21633];
                
                r_data[21635] <= r_data[21634];
                
                r_data[21636] <= r_data[21635];
                
                r_data[21637] <= r_data[21636];
                
                r_data[21638] <= r_data[21637];
                
                r_data[21639] <= r_data[21638];
                
                r_data[21640] <= r_data[21639];
                
                r_data[21641] <= r_data[21640];
                
                r_data[21642] <= r_data[21641];
                
                r_data[21643] <= r_data[21642];
                
                r_data[21644] <= r_data[21643];
                
                r_data[21645] <= r_data[21644];
                
                r_data[21646] <= r_data[21645];
                
                r_data[21647] <= r_data[21646];
                
                r_data[21648] <= r_data[21647];
                
                r_data[21649] <= r_data[21648];
                
                r_data[21650] <= r_data[21649];
                
                r_data[21651] <= r_data[21650];
                
                r_data[21652] <= r_data[21651];
                
                r_data[21653] <= r_data[21652];
                
                r_data[21654] <= r_data[21653];
                
                r_data[21655] <= r_data[21654];
                
                r_data[21656] <= r_data[21655];
                
                r_data[21657] <= r_data[21656];
                
                r_data[21658] <= r_data[21657];
                
                r_data[21659] <= r_data[21658];
                
                r_data[21660] <= r_data[21659];
                
                r_data[21661] <= r_data[21660];
                
                r_data[21662] <= r_data[21661];
                
                r_data[21663] <= r_data[21662];
                
                r_data[21664] <= r_data[21663];
                
                r_data[21665] <= r_data[21664];
                
                r_data[21666] <= r_data[21665];
                
                r_data[21667] <= r_data[21666];
                
                r_data[21668] <= r_data[21667];
                
                r_data[21669] <= r_data[21668];
                
                r_data[21670] <= r_data[21669];
                
                r_data[21671] <= r_data[21670];
                
                r_data[21672] <= r_data[21671];
                
                r_data[21673] <= r_data[21672];
                
                r_data[21674] <= r_data[21673];
                
                r_data[21675] <= r_data[21674];
                
                r_data[21676] <= r_data[21675];
                
                r_data[21677] <= r_data[21676];
                
                r_data[21678] <= r_data[21677];
                
                r_data[21679] <= r_data[21678];
                
                r_data[21680] <= r_data[21679];
                
                r_data[21681] <= r_data[21680];
                
                r_data[21682] <= r_data[21681];
                
                r_data[21683] <= r_data[21682];
                
                r_data[21684] <= r_data[21683];
                
                r_data[21685] <= r_data[21684];
                
                r_data[21686] <= r_data[21685];
                
                r_data[21687] <= r_data[21686];
                
                r_data[21688] <= r_data[21687];
                
                r_data[21689] <= r_data[21688];
                
                r_data[21690] <= r_data[21689];
                
                r_data[21691] <= r_data[21690];
                
                r_data[21692] <= r_data[21691];
                
                r_data[21693] <= r_data[21692];
                
                r_data[21694] <= r_data[21693];
                
                r_data[21695] <= r_data[21694];
                
                r_data[21696] <= r_data[21695];
                
                r_data[21697] <= r_data[21696];
                
                r_data[21698] <= r_data[21697];
                
                r_data[21699] <= r_data[21698];
                
                r_data[21700] <= r_data[21699];
                
                r_data[21701] <= r_data[21700];
                
                r_data[21702] <= r_data[21701];
                
                r_data[21703] <= r_data[21702];
                
                r_data[21704] <= r_data[21703];
                
                r_data[21705] <= r_data[21704];
                
                r_data[21706] <= r_data[21705];
                
                r_data[21707] <= r_data[21706];
                
                r_data[21708] <= r_data[21707];
                
                r_data[21709] <= r_data[21708];
                
                r_data[21710] <= r_data[21709];
                
                r_data[21711] <= r_data[21710];
                
                r_data[21712] <= r_data[21711];
                
                r_data[21713] <= r_data[21712];
                
                r_data[21714] <= r_data[21713];
                
                r_data[21715] <= r_data[21714];
                
                r_data[21716] <= r_data[21715];
                
                r_data[21717] <= r_data[21716];
                
                r_data[21718] <= r_data[21717];
                
                r_data[21719] <= r_data[21718];
                
                r_data[21720] <= r_data[21719];
                
                r_data[21721] <= r_data[21720];
                
                r_data[21722] <= r_data[21721];
                
                r_data[21723] <= r_data[21722];
                
                r_data[21724] <= r_data[21723];
                
                r_data[21725] <= r_data[21724];
                
                r_data[21726] <= r_data[21725];
                
                r_data[21727] <= r_data[21726];
                
                r_data[21728] <= r_data[21727];
                
                r_data[21729] <= r_data[21728];
                
                r_data[21730] <= r_data[21729];
                
                r_data[21731] <= r_data[21730];
                
                r_data[21732] <= r_data[21731];
                
                r_data[21733] <= r_data[21732];
                
                r_data[21734] <= r_data[21733];
                
                r_data[21735] <= r_data[21734];
                
                r_data[21736] <= r_data[21735];
                
                r_data[21737] <= r_data[21736];
                
                r_data[21738] <= r_data[21737];
                
                r_data[21739] <= r_data[21738];
                
                r_data[21740] <= r_data[21739];
                
                r_data[21741] <= r_data[21740];
                
                r_data[21742] <= r_data[21741];
                
                r_data[21743] <= r_data[21742];
                
                r_data[21744] <= r_data[21743];
                
                r_data[21745] <= r_data[21744];
                
                r_data[21746] <= r_data[21745];
                
                r_data[21747] <= r_data[21746];
                
                r_data[21748] <= r_data[21747];
                
                r_data[21749] <= r_data[21748];
                
                r_data[21750] <= r_data[21749];
                
                r_data[21751] <= r_data[21750];
                
                r_data[21752] <= r_data[21751];
                
                r_data[21753] <= r_data[21752];
                
                r_data[21754] <= r_data[21753];
                
                r_data[21755] <= r_data[21754];
                
                r_data[21756] <= r_data[21755];
                
                r_data[21757] <= r_data[21756];
                
                r_data[21758] <= r_data[21757];
                
                r_data[21759] <= r_data[21758];
                
                r_data[21760] <= r_data[21759];
                
                r_data[21761] <= r_data[21760];
                
                r_data[21762] <= r_data[21761];
                
                r_data[21763] <= r_data[21762];
                
                r_data[21764] <= r_data[21763];
                
                r_data[21765] <= r_data[21764];
                
                r_data[21766] <= r_data[21765];
                
                r_data[21767] <= r_data[21766];
                
                r_data[21768] <= r_data[21767];
                
                r_data[21769] <= r_data[21768];
                
                r_data[21770] <= r_data[21769];
                
                r_data[21771] <= r_data[21770];
                
                r_data[21772] <= r_data[21771];
                
                r_data[21773] <= r_data[21772];
                
                r_data[21774] <= r_data[21773];
                
                r_data[21775] <= r_data[21774];
                
                r_data[21776] <= r_data[21775];
                
                r_data[21777] <= r_data[21776];
                
                r_data[21778] <= r_data[21777];
                
                r_data[21779] <= r_data[21778];
                
                r_data[21780] <= r_data[21779];
                
                r_data[21781] <= r_data[21780];
                
                r_data[21782] <= r_data[21781];
                
                r_data[21783] <= r_data[21782];
                
                r_data[21784] <= r_data[21783];
                
                r_data[21785] <= r_data[21784];
                
                r_data[21786] <= r_data[21785];
                
                r_data[21787] <= r_data[21786];
                
                r_data[21788] <= r_data[21787];
                
                r_data[21789] <= r_data[21788];
                
                r_data[21790] <= r_data[21789];
                
                r_data[21791] <= r_data[21790];
                
                r_data[21792] <= r_data[21791];
                
                r_data[21793] <= r_data[21792];
                
                r_data[21794] <= r_data[21793];
                
                r_data[21795] <= r_data[21794];
                
                r_data[21796] <= r_data[21795];
                
                r_data[21797] <= r_data[21796];
                
                r_data[21798] <= r_data[21797];
                
                r_data[21799] <= r_data[21798];
                
                r_data[21800] <= r_data[21799];
                
                r_data[21801] <= r_data[21800];
                
                r_data[21802] <= r_data[21801];
                
                r_data[21803] <= r_data[21802];
                
                r_data[21804] <= r_data[21803];
                
                r_data[21805] <= r_data[21804];
                
                r_data[21806] <= r_data[21805];
                
                r_data[21807] <= r_data[21806];
                
                r_data[21808] <= r_data[21807];
                
                r_data[21809] <= r_data[21808];
                
                r_data[21810] <= r_data[21809];
                
                r_data[21811] <= r_data[21810];
                
                r_data[21812] <= r_data[21811];
                
                r_data[21813] <= r_data[21812];
                
                r_data[21814] <= r_data[21813];
                
                r_data[21815] <= r_data[21814];
                
                r_data[21816] <= r_data[21815];
                
                r_data[21817] <= r_data[21816];
                
                r_data[21818] <= r_data[21817];
                
                r_data[21819] <= r_data[21818];
                
                r_data[21820] <= r_data[21819];
                
                r_data[21821] <= r_data[21820];
                
                r_data[21822] <= r_data[21821];
                
                r_data[21823] <= r_data[21822];
                
                r_data[21824] <= r_data[21823];
                
                r_data[21825] <= r_data[21824];
                
                r_data[21826] <= r_data[21825];
                
                r_data[21827] <= r_data[21826];
                
                r_data[21828] <= r_data[21827];
                
                r_data[21829] <= r_data[21828];
                
                r_data[21830] <= r_data[21829];
                
                r_data[21831] <= r_data[21830];
                
                r_data[21832] <= r_data[21831];
                
                r_data[21833] <= r_data[21832];
                
                r_data[21834] <= r_data[21833];
                
                r_data[21835] <= r_data[21834];
                
                r_data[21836] <= r_data[21835];
                
                r_data[21837] <= r_data[21836];
                
                r_data[21838] <= r_data[21837];
                
                r_data[21839] <= r_data[21838];
                
                r_data[21840] <= r_data[21839];
                
                r_data[21841] <= r_data[21840];
                
                r_data[21842] <= r_data[21841];
                
                r_data[21843] <= r_data[21842];
                
                r_data[21844] <= r_data[21843];
                
                r_data[21845] <= r_data[21844];
                
                r_data[21846] <= r_data[21845];
                
                r_data[21847] <= r_data[21846];
                
                r_data[21848] <= r_data[21847];
                
                r_data[21849] <= r_data[21848];
                
                r_data[21850] <= r_data[21849];
                
                r_data[21851] <= r_data[21850];
                
                r_data[21852] <= r_data[21851];
                
                r_data[21853] <= r_data[21852];
                
                r_data[21854] <= r_data[21853];
                
                r_data[21855] <= r_data[21854];
                
                r_data[21856] <= r_data[21855];
                
                r_data[21857] <= r_data[21856];
                
                r_data[21858] <= r_data[21857];
                
                r_data[21859] <= r_data[21858];
                
                r_data[21860] <= r_data[21859];
                
                r_data[21861] <= r_data[21860];
                
                r_data[21862] <= r_data[21861];
                
                r_data[21863] <= r_data[21862];
                
                r_data[21864] <= r_data[21863];
                
                r_data[21865] <= r_data[21864];
                
                r_data[21866] <= r_data[21865];
                
                r_data[21867] <= r_data[21866];
                
                r_data[21868] <= r_data[21867];
                
                r_data[21869] <= r_data[21868];
                
                r_data[21870] <= r_data[21869];
                
                r_data[21871] <= r_data[21870];
                
                r_data[21872] <= r_data[21871];
                
                r_data[21873] <= r_data[21872];
                
                r_data[21874] <= r_data[21873];
                
                r_data[21875] <= r_data[21874];
                
                r_data[21876] <= r_data[21875];
                
                r_data[21877] <= r_data[21876];
                
                r_data[21878] <= r_data[21877];
                
                r_data[21879] <= r_data[21878];
                
                r_data[21880] <= r_data[21879];
                
                r_data[21881] <= r_data[21880];
                
                r_data[21882] <= r_data[21881];
                
                r_data[21883] <= r_data[21882];
                
                r_data[21884] <= r_data[21883];
                
                r_data[21885] <= r_data[21884];
                
                r_data[21886] <= r_data[21885];
                
                r_data[21887] <= r_data[21886];
                
                r_data[21888] <= r_data[21887];
                
                r_data[21889] <= r_data[21888];
                
                r_data[21890] <= r_data[21889];
                
                r_data[21891] <= r_data[21890];
                
                r_data[21892] <= r_data[21891];
                
                r_data[21893] <= r_data[21892];
                
                r_data[21894] <= r_data[21893];
                
                r_data[21895] <= r_data[21894];
                
                r_data[21896] <= r_data[21895];
                
                r_data[21897] <= r_data[21896];
                
                r_data[21898] <= r_data[21897];
                
                r_data[21899] <= r_data[21898];
                
                r_data[21900] <= r_data[21899];
                
                r_data[21901] <= r_data[21900];
                
                r_data[21902] <= r_data[21901];
                
                r_data[21903] <= r_data[21902];
                
                r_data[21904] <= r_data[21903];
                
                r_data[21905] <= r_data[21904];
                
                r_data[21906] <= r_data[21905];
                
                r_data[21907] <= r_data[21906];
                
                r_data[21908] <= r_data[21907];
                
                r_data[21909] <= r_data[21908];
                
                r_data[21910] <= r_data[21909];
                
                r_data[21911] <= r_data[21910];
                
                r_data[21912] <= r_data[21911];
                
                r_data[21913] <= r_data[21912];
                
                r_data[21914] <= r_data[21913];
                
                r_data[21915] <= r_data[21914];
                
                r_data[21916] <= r_data[21915];
                
                r_data[21917] <= r_data[21916];
                
                r_data[21918] <= r_data[21917];
                
                r_data[21919] <= r_data[21918];
                
                r_data[21920] <= r_data[21919];
                
                r_data[21921] <= r_data[21920];
                
                r_data[21922] <= r_data[21921];
                
                r_data[21923] <= r_data[21922];
                
                r_data[21924] <= r_data[21923];
                
                r_data[21925] <= r_data[21924];
                
                r_data[21926] <= r_data[21925];
                
                r_data[21927] <= r_data[21926];
                
                r_data[21928] <= r_data[21927];
                
                r_data[21929] <= r_data[21928];
                
                r_data[21930] <= r_data[21929];
                
                r_data[21931] <= r_data[21930];
                
                r_data[21932] <= r_data[21931];
                
                r_data[21933] <= r_data[21932];
                
                r_data[21934] <= r_data[21933];
                
                r_data[21935] <= r_data[21934];
                
                r_data[21936] <= r_data[21935];
                
                r_data[21937] <= r_data[21936];
                
                r_data[21938] <= r_data[21937];
                
                r_data[21939] <= r_data[21938];
                
                r_data[21940] <= r_data[21939];
                
                r_data[21941] <= r_data[21940];
                
                r_data[21942] <= r_data[21941];
                
                r_data[21943] <= r_data[21942];
                
                r_data[21944] <= r_data[21943];
                
                r_data[21945] <= r_data[21944];
                
                r_data[21946] <= r_data[21945];
                
                r_data[21947] <= r_data[21946];
                
                r_data[21948] <= r_data[21947];
                
                r_data[21949] <= r_data[21948];
                
                r_data[21950] <= r_data[21949];
                
                r_data[21951] <= r_data[21950];
                
                r_data[21952] <= r_data[21951];
                
                r_data[21953] <= r_data[21952];
                
                r_data[21954] <= r_data[21953];
                
                r_data[21955] <= r_data[21954];
                
                r_data[21956] <= r_data[21955];
                
                r_data[21957] <= r_data[21956];
                
                r_data[21958] <= r_data[21957];
                
                r_data[21959] <= r_data[21958];
                
                r_data[21960] <= r_data[21959];
                
                r_data[21961] <= r_data[21960];
                
                r_data[21962] <= r_data[21961];
                
                r_data[21963] <= r_data[21962];
                
                r_data[21964] <= r_data[21963];
                
                r_data[21965] <= r_data[21964];
                
                r_data[21966] <= r_data[21965];
                
                r_data[21967] <= r_data[21966];
                
                r_data[21968] <= r_data[21967];
                
                r_data[21969] <= r_data[21968];
                
                r_data[21970] <= r_data[21969];
                
                r_data[21971] <= r_data[21970];
                
                r_data[21972] <= r_data[21971];
                
                r_data[21973] <= r_data[21972];
                
                r_data[21974] <= r_data[21973];
                
                r_data[21975] <= r_data[21974];
                
                r_data[21976] <= r_data[21975];
                
                r_data[21977] <= r_data[21976];
                
                r_data[21978] <= r_data[21977];
                
                r_data[21979] <= r_data[21978];
                
                r_data[21980] <= r_data[21979];
                
                r_data[21981] <= r_data[21980];
                
                r_data[21982] <= r_data[21981];
                
                r_data[21983] <= r_data[21982];
                
                r_data[21984] <= r_data[21983];
                
                r_data[21985] <= r_data[21984];
                
                r_data[21986] <= r_data[21985];
                
                r_data[21987] <= r_data[21986];
                
                r_data[21988] <= r_data[21987];
                
                r_data[21989] <= r_data[21988];
                
                r_data[21990] <= r_data[21989];
                
                r_data[21991] <= r_data[21990];
                
                r_data[21992] <= r_data[21991];
                
                r_data[21993] <= r_data[21992];
                
                r_data[21994] <= r_data[21993];
                
                r_data[21995] <= r_data[21994];
                
                r_data[21996] <= r_data[21995];
                
                r_data[21997] <= r_data[21996];
                
                r_data[21998] <= r_data[21997];
                
                r_data[21999] <= r_data[21998];
                
                r_data[22000] <= r_data[21999];
                
                r_data[22001] <= r_data[22000];
                
                r_data[22002] <= r_data[22001];
                
                r_data[22003] <= r_data[22002];
                
                r_data[22004] <= r_data[22003];
                
                r_data[22005] <= r_data[22004];
                
                r_data[22006] <= r_data[22005];
                
                r_data[22007] <= r_data[22006];
                
                r_data[22008] <= r_data[22007];
                
                r_data[22009] <= r_data[22008];
                
                r_data[22010] <= r_data[22009];
                
                r_data[22011] <= r_data[22010];
                
                r_data[22012] <= r_data[22011];
                
                r_data[22013] <= r_data[22012];
                
                r_data[22014] <= r_data[22013];
                
                r_data[22015] <= r_data[22014];
                
                r_data[22016] <= r_data[22015];
                
                r_data[22017] <= r_data[22016];
                
                r_data[22018] <= r_data[22017];
                
                r_data[22019] <= r_data[22018];
                
                r_data[22020] <= r_data[22019];
                
                r_data[22021] <= r_data[22020];
                
                r_data[22022] <= r_data[22021];
                
                r_data[22023] <= r_data[22022];
                
                r_data[22024] <= r_data[22023];
                
                r_data[22025] <= r_data[22024];
                
                r_data[22026] <= r_data[22025];
                
                r_data[22027] <= r_data[22026];
                
                r_data[22028] <= r_data[22027];
                
                r_data[22029] <= r_data[22028];
                
                r_data[22030] <= r_data[22029];
                
                r_data[22031] <= r_data[22030];
                
                r_data[22032] <= r_data[22031];
                
                r_data[22033] <= r_data[22032];
                
                r_data[22034] <= r_data[22033];
                
                r_data[22035] <= r_data[22034];
                
                r_data[22036] <= r_data[22035];
                
                r_data[22037] <= r_data[22036];
                
                r_data[22038] <= r_data[22037];
                
                r_data[22039] <= r_data[22038];
                
                r_data[22040] <= r_data[22039];
                
                r_data[22041] <= r_data[22040];
                
                r_data[22042] <= r_data[22041];
                
                r_data[22043] <= r_data[22042];
                
                r_data[22044] <= r_data[22043];
                
                r_data[22045] <= r_data[22044];
                
                r_data[22046] <= r_data[22045];
                
                r_data[22047] <= r_data[22046];
                
                r_data[22048] <= r_data[22047];
                
                r_data[22049] <= r_data[22048];
                
                r_data[22050] <= r_data[22049];
                
                r_data[22051] <= r_data[22050];
                
                r_data[22052] <= r_data[22051];
                
                r_data[22053] <= r_data[22052];
                
                r_data[22054] <= r_data[22053];
                
                r_data[22055] <= r_data[22054];
                
                r_data[22056] <= r_data[22055];
                
                r_data[22057] <= r_data[22056];
                
                r_data[22058] <= r_data[22057];
                
                r_data[22059] <= r_data[22058];
                
                r_data[22060] <= r_data[22059];
                
                r_data[22061] <= r_data[22060];
                
                r_data[22062] <= r_data[22061];
                
                r_data[22063] <= r_data[22062];
                
                r_data[22064] <= r_data[22063];
                
                r_data[22065] <= r_data[22064];
                
                r_data[22066] <= r_data[22065];
                
                r_data[22067] <= r_data[22066];
                
                r_data[22068] <= r_data[22067];
                
                r_data[22069] <= r_data[22068];
                
                r_data[22070] <= r_data[22069];
                
                r_data[22071] <= r_data[22070];
                
                r_data[22072] <= r_data[22071];
                
                r_data[22073] <= r_data[22072];
                
                r_data[22074] <= r_data[22073];
                
                r_data[22075] <= r_data[22074];
                
                r_data[22076] <= r_data[22075];
                
                r_data[22077] <= r_data[22076];
                
                r_data[22078] <= r_data[22077];
                
                r_data[22079] <= r_data[22078];
                
                r_data[22080] <= r_data[22079];
                
                r_data[22081] <= r_data[22080];
                
                r_data[22082] <= r_data[22081];
                
                r_data[22083] <= r_data[22082];
                
                r_data[22084] <= r_data[22083];
                
                r_data[22085] <= r_data[22084];
                
                r_data[22086] <= r_data[22085];
                
                r_data[22087] <= r_data[22086];
                
                r_data[22088] <= r_data[22087];
                
                r_data[22089] <= r_data[22088];
                
                r_data[22090] <= r_data[22089];
                
                r_data[22091] <= r_data[22090];
                
                r_data[22092] <= r_data[22091];
                
                r_data[22093] <= r_data[22092];
                
                r_data[22094] <= r_data[22093];
                
                r_data[22095] <= r_data[22094];
                
                r_data[22096] <= r_data[22095];
                
                r_data[22097] <= r_data[22096];
                
                r_data[22098] <= r_data[22097];
                
                r_data[22099] <= r_data[22098];
                
                r_data[22100] <= r_data[22099];
                
                r_data[22101] <= r_data[22100];
                
                r_data[22102] <= r_data[22101];
                
                r_data[22103] <= r_data[22102];
                
                r_data[22104] <= r_data[22103];
                
                r_data[22105] <= r_data[22104];
                
                r_data[22106] <= r_data[22105];
                
                r_data[22107] <= r_data[22106];
                
                r_data[22108] <= r_data[22107];
                
                r_data[22109] <= r_data[22108];
                
                r_data[22110] <= r_data[22109];
                
                r_data[22111] <= r_data[22110];
                
                r_data[22112] <= r_data[22111];
                
                r_data[22113] <= r_data[22112];
                
                r_data[22114] <= r_data[22113];
                
                r_data[22115] <= r_data[22114];
                
                r_data[22116] <= r_data[22115];
                
                r_data[22117] <= r_data[22116];
                
                r_data[22118] <= r_data[22117];
                
                r_data[22119] <= r_data[22118];
                
                r_data[22120] <= r_data[22119];
                
                r_data[22121] <= r_data[22120];
                
                r_data[22122] <= r_data[22121];
                
                r_data[22123] <= r_data[22122];
                
                r_data[22124] <= r_data[22123];
                
                r_data[22125] <= r_data[22124];
                
                r_data[22126] <= r_data[22125];
                
                r_data[22127] <= r_data[22126];
                
                r_data[22128] <= r_data[22127];
                
                r_data[22129] <= r_data[22128];
                
                r_data[22130] <= r_data[22129];
                
                r_data[22131] <= r_data[22130];
                
                r_data[22132] <= r_data[22131];
                
                r_data[22133] <= r_data[22132];
                
                r_data[22134] <= r_data[22133];
                
                r_data[22135] <= r_data[22134];
                
                r_data[22136] <= r_data[22135];
                
                r_data[22137] <= r_data[22136];
                
                r_data[22138] <= r_data[22137];
                
                r_data[22139] <= r_data[22138];
                
                r_data[22140] <= r_data[22139];
                
                r_data[22141] <= r_data[22140];
                
                r_data[22142] <= r_data[22141];
                
                r_data[22143] <= r_data[22142];
                
                r_data[22144] <= r_data[22143];
                
                r_data[22145] <= r_data[22144];
                
                r_data[22146] <= r_data[22145];
                
                r_data[22147] <= r_data[22146];
                
                r_data[22148] <= r_data[22147];
                
                r_data[22149] <= r_data[22148];
                
                r_data[22150] <= r_data[22149];
                
                r_data[22151] <= r_data[22150];
                
                r_data[22152] <= r_data[22151];
                
                r_data[22153] <= r_data[22152];
                
                r_data[22154] <= r_data[22153];
                
                r_data[22155] <= r_data[22154];
                
                r_data[22156] <= r_data[22155];
                
                r_data[22157] <= r_data[22156];
                
                r_data[22158] <= r_data[22157];
                
                r_data[22159] <= r_data[22158];
                
                r_data[22160] <= r_data[22159];
                
                r_data[22161] <= r_data[22160];
                
                r_data[22162] <= r_data[22161];
                
                r_data[22163] <= r_data[22162];
                
                r_data[22164] <= r_data[22163];
                
                r_data[22165] <= r_data[22164];
                
                r_data[22166] <= r_data[22165];
                
                r_data[22167] <= r_data[22166];
                
                r_data[22168] <= r_data[22167];
                
                r_data[22169] <= r_data[22168];
                
                r_data[22170] <= r_data[22169];
                
                r_data[22171] <= r_data[22170];
                
                r_data[22172] <= r_data[22171];
                
                r_data[22173] <= r_data[22172];
                
                r_data[22174] <= r_data[22173];
                
                r_data[22175] <= r_data[22174];
                
                r_data[22176] <= r_data[22175];
                
                r_data[22177] <= r_data[22176];
                
                r_data[22178] <= r_data[22177];
                
                r_data[22179] <= r_data[22178];
                
                r_data[22180] <= r_data[22179];
                
                r_data[22181] <= r_data[22180];
                
                r_data[22182] <= r_data[22181];
                
                r_data[22183] <= r_data[22182];
                
                r_data[22184] <= r_data[22183];
                
                r_data[22185] <= r_data[22184];
                
                r_data[22186] <= r_data[22185];
                
                r_data[22187] <= r_data[22186];
                
                r_data[22188] <= r_data[22187];
                
                r_data[22189] <= r_data[22188];
                
                r_data[22190] <= r_data[22189];
                
                r_data[22191] <= r_data[22190];
                
                r_data[22192] <= r_data[22191];
                
                r_data[22193] <= r_data[22192];
                
                r_data[22194] <= r_data[22193];
                
                r_data[22195] <= r_data[22194];
                
                r_data[22196] <= r_data[22195];
                
                r_data[22197] <= r_data[22196];
                
                r_data[22198] <= r_data[22197];
                
                r_data[22199] <= r_data[22198];
                
                r_data[22200] <= r_data[22199];
                
                r_data[22201] <= r_data[22200];
                
                r_data[22202] <= r_data[22201];
                
                r_data[22203] <= r_data[22202];
                
                r_data[22204] <= r_data[22203];
                
                r_data[22205] <= r_data[22204];
                
                r_data[22206] <= r_data[22205];
                
                r_data[22207] <= r_data[22206];
                
                r_data[22208] <= r_data[22207];
                
                r_data[22209] <= r_data[22208];
                
                r_data[22210] <= r_data[22209];
                
                r_data[22211] <= r_data[22210];
                
                r_data[22212] <= r_data[22211];
                
                r_data[22213] <= r_data[22212];
                
                r_data[22214] <= r_data[22213];
                
                r_data[22215] <= r_data[22214];
                
                r_data[22216] <= r_data[22215];
                
                r_data[22217] <= r_data[22216];
                
                r_data[22218] <= r_data[22217];
                
                r_data[22219] <= r_data[22218];
                
                r_data[22220] <= r_data[22219];
                
                r_data[22221] <= r_data[22220];
                
                r_data[22222] <= r_data[22221];
                
                r_data[22223] <= r_data[22222];
                
                r_data[22224] <= r_data[22223];
                
                r_data[22225] <= r_data[22224];
                
                r_data[22226] <= r_data[22225];
                
                r_data[22227] <= r_data[22226];
                
                r_data[22228] <= r_data[22227];
                
                r_data[22229] <= r_data[22228];
                
                r_data[22230] <= r_data[22229];
                
                r_data[22231] <= r_data[22230];
                
                r_data[22232] <= r_data[22231];
                
                r_data[22233] <= r_data[22232];
                
                r_data[22234] <= r_data[22233];
                
                r_data[22235] <= r_data[22234];
                
                r_data[22236] <= r_data[22235];
                
                r_data[22237] <= r_data[22236];
                
                r_data[22238] <= r_data[22237];
                
                r_data[22239] <= r_data[22238];
                
                r_data[22240] <= r_data[22239];
                
                r_data[22241] <= r_data[22240];
                
                r_data[22242] <= r_data[22241];
                
                r_data[22243] <= r_data[22242];
                
                r_data[22244] <= r_data[22243];
                
                r_data[22245] <= r_data[22244];
                
                r_data[22246] <= r_data[22245];
                
                r_data[22247] <= r_data[22246];
                
                r_data[22248] <= r_data[22247];
                
                r_data[22249] <= r_data[22248];
                
                r_data[22250] <= r_data[22249];
                
                r_data[22251] <= r_data[22250];
                
                r_data[22252] <= r_data[22251];
                
                r_data[22253] <= r_data[22252];
                
                r_data[22254] <= r_data[22253];
                
                r_data[22255] <= r_data[22254];
                
                r_data[22256] <= r_data[22255];
                
                r_data[22257] <= r_data[22256];
                
                r_data[22258] <= r_data[22257];
                
                r_data[22259] <= r_data[22258];
                
                r_data[22260] <= r_data[22259];
                
                r_data[22261] <= r_data[22260];
                
                r_data[22262] <= r_data[22261];
                
                r_data[22263] <= r_data[22262];
                
                r_data[22264] <= r_data[22263];
                
                r_data[22265] <= r_data[22264];
                
                r_data[22266] <= r_data[22265];
                
                r_data[22267] <= r_data[22266];
                
                r_data[22268] <= r_data[22267];
                
                r_data[22269] <= r_data[22268];
                
                r_data[22270] <= r_data[22269];
                
                r_data[22271] <= r_data[22270];
                
                r_data[22272] <= r_data[22271];
                
                r_data[22273] <= r_data[22272];
                
                r_data[22274] <= r_data[22273];
                
                r_data[22275] <= r_data[22274];
                
                r_data[22276] <= r_data[22275];
                
                r_data[22277] <= r_data[22276];
                
                r_data[22278] <= r_data[22277];
                
                r_data[22279] <= r_data[22278];
                
                r_data[22280] <= r_data[22279];
                
                r_data[22281] <= r_data[22280];
                
                r_data[22282] <= r_data[22281];
                
                r_data[22283] <= r_data[22282];
                
                r_data[22284] <= r_data[22283];
                
                r_data[22285] <= r_data[22284];
                
                r_data[22286] <= r_data[22285];
                
                r_data[22287] <= r_data[22286];
                
                r_data[22288] <= r_data[22287];
                
                r_data[22289] <= r_data[22288];
                
                r_data[22290] <= r_data[22289];
                
                r_data[22291] <= r_data[22290];
                
                r_data[22292] <= r_data[22291];
                
                r_data[22293] <= r_data[22292];
                
                r_data[22294] <= r_data[22293];
                
                r_data[22295] <= r_data[22294];
                
                r_data[22296] <= r_data[22295];
                
                r_data[22297] <= r_data[22296];
                
                r_data[22298] <= r_data[22297];
                
                r_data[22299] <= r_data[22298];
                
                r_data[22300] <= r_data[22299];
                
                r_data[22301] <= r_data[22300];
                
                r_data[22302] <= r_data[22301];
                
                r_data[22303] <= r_data[22302];
                
                r_data[22304] <= r_data[22303];
                
                r_data[22305] <= r_data[22304];
                
                r_data[22306] <= r_data[22305];
                
                r_data[22307] <= r_data[22306];
                
                r_data[22308] <= r_data[22307];
                
                r_data[22309] <= r_data[22308];
                
                r_data[22310] <= r_data[22309];
                
                r_data[22311] <= r_data[22310];
                
                r_data[22312] <= r_data[22311];
                
                r_data[22313] <= r_data[22312];
                
                r_data[22314] <= r_data[22313];
                
                r_data[22315] <= r_data[22314];
                
                r_data[22316] <= r_data[22315];
                
                r_data[22317] <= r_data[22316];
                
                r_data[22318] <= r_data[22317];
                
                r_data[22319] <= r_data[22318];
                
                r_data[22320] <= r_data[22319];
                
                r_data[22321] <= r_data[22320];
                
                r_data[22322] <= r_data[22321];
                
                r_data[22323] <= r_data[22322];
                
                r_data[22324] <= r_data[22323];
                
                r_data[22325] <= r_data[22324];
                
                r_data[22326] <= r_data[22325];
                
                r_data[22327] <= r_data[22326];
                
                r_data[22328] <= r_data[22327];
                
                r_data[22329] <= r_data[22328];
                
                r_data[22330] <= r_data[22329];
                
                r_data[22331] <= r_data[22330];
                
                r_data[22332] <= r_data[22331];
                
                r_data[22333] <= r_data[22332];
                
                r_data[22334] <= r_data[22333];
                
                r_data[22335] <= r_data[22334];
                
                r_data[22336] <= r_data[22335];
                
                r_data[22337] <= r_data[22336];
                
                r_data[22338] <= r_data[22337];
                
                r_data[22339] <= r_data[22338];
                
                r_data[22340] <= r_data[22339];
                
                r_data[22341] <= r_data[22340];
                
                r_data[22342] <= r_data[22341];
                
                r_data[22343] <= r_data[22342];
                
                r_data[22344] <= r_data[22343];
                
                r_data[22345] <= r_data[22344];
                
                r_data[22346] <= r_data[22345];
                
                r_data[22347] <= r_data[22346];
                
                r_data[22348] <= r_data[22347];
                
                r_data[22349] <= r_data[22348];
                
                r_data[22350] <= r_data[22349];
                
                r_data[22351] <= r_data[22350];
                
                r_data[22352] <= r_data[22351];
                
                r_data[22353] <= r_data[22352];
                
                r_data[22354] <= r_data[22353];
                
                r_data[22355] <= r_data[22354];
                
                r_data[22356] <= r_data[22355];
                
                r_data[22357] <= r_data[22356];
                
                r_data[22358] <= r_data[22357];
                
                r_data[22359] <= r_data[22358];
                
                r_data[22360] <= r_data[22359];
                
                r_data[22361] <= r_data[22360];
                
                r_data[22362] <= r_data[22361];
                
                r_data[22363] <= r_data[22362];
                
                r_data[22364] <= r_data[22363];
                
                r_data[22365] <= r_data[22364];
                
                r_data[22366] <= r_data[22365];
                
                r_data[22367] <= r_data[22366];
                
                r_data[22368] <= r_data[22367];
                
                r_data[22369] <= r_data[22368];
                
                r_data[22370] <= r_data[22369];
                
                r_data[22371] <= r_data[22370];
                
                r_data[22372] <= r_data[22371];
                
                r_data[22373] <= r_data[22372];
                
                r_data[22374] <= r_data[22373];
                
                r_data[22375] <= r_data[22374];
                
                r_data[22376] <= r_data[22375];
                
                r_data[22377] <= r_data[22376];
                
                r_data[22378] <= r_data[22377];
                
                r_data[22379] <= r_data[22378];
                
                r_data[22380] <= r_data[22379];
                
                r_data[22381] <= r_data[22380];
                
                r_data[22382] <= r_data[22381];
                
                r_data[22383] <= r_data[22382];
                
                r_data[22384] <= r_data[22383];
                
                r_data[22385] <= r_data[22384];
                
                r_data[22386] <= r_data[22385];
                
                r_data[22387] <= r_data[22386];
                
                r_data[22388] <= r_data[22387];
                
                r_data[22389] <= r_data[22388];
                
                r_data[22390] <= r_data[22389];
                
                r_data[22391] <= r_data[22390];
                
                r_data[22392] <= r_data[22391];
                
                r_data[22393] <= r_data[22392];
                
                r_data[22394] <= r_data[22393];
                
                r_data[22395] <= r_data[22394];
                
                r_data[22396] <= r_data[22395];
                
                r_data[22397] <= r_data[22396];
                
                r_data[22398] <= r_data[22397];
                
                r_data[22399] <= r_data[22398];
                
                r_data[22400] <= r_data[22399];
                
                r_data[22401] <= r_data[22400];
                
                r_data[22402] <= r_data[22401];
                
                r_data[22403] <= r_data[22402];
                
                r_data[22404] <= r_data[22403];
                
                r_data[22405] <= r_data[22404];
                
                r_data[22406] <= r_data[22405];
                
                r_data[22407] <= r_data[22406];
                
                r_data[22408] <= r_data[22407];
                
                r_data[22409] <= r_data[22408];
                
                r_data[22410] <= r_data[22409];
                
                r_data[22411] <= r_data[22410];
                
                r_data[22412] <= r_data[22411];
                
                r_data[22413] <= r_data[22412];
                
                r_data[22414] <= r_data[22413];
                
                r_data[22415] <= r_data[22414];
                
                r_data[22416] <= r_data[22415];
                
                r_data[22417] <= r_data[22416];
                
                r_data[22418] <= r_data[22417];
                
                r_data[22419] <= r_data[22418];
                
                r_data[22420] <= r_data[22419];
                
                r_data[22421] <= r_data[22420];
                
                r_data[22422] <= r_data[22421];
                
                r_data[22423] <= r_data[22422];
                
                r_data[22424] <= r_data[22423];
                
                r_data[22425] <= r_data[22424];
                
                r_data[22426] <= r_data[22425];
                
                r_data[22427] <= r_data[22426];
                
                r_data[22428] <= r_data[22427];
                
                r_data[22429] <= r_data[22428];
                
                r_data[22430] <= r_data[22429];
                
                r_data[22431] <= r_data[22430];
                
                r_data[22432] <= r_data[22431];
                
                r_data[22433] <= r_data[22432];
                
                r_data[22434] <= r_data[22433];
                
                r_data[22435] <= r_data[22434];
                
                r_data[22436] <= r_data[22435];
                
                r_data[22437] <= r_data[22436];
                
                r_data[22438] <= r_data[22437];
                
                r_data[22439] <= r_data[22438];
                
                r_data[22440] <= r_data[22439];
                
                r_data[22441] <= r_data[22440];
                
                r_data[22442] <= r_data[22441];
                
                r_data[22443] <= r_data[22442];
                
                r_data[22444] <= r_data[22443];
                
                r_data[22445] <= r_data[22444];
                
                r_data[22446] <= r_data[22445];
                
                r_data[22447] <= r_data[22446];
                
                r_data[22448] <= r_data[22447];
                
                r_data[22449] <= r_data[22448];
                
                r_data[22450] <= r_data[22449];
                
                r_data[22451] <= r_data[22450];
                
                r_data[22452] <= r_data[22451];
                
                r_data[22453] <= r_data[22452];
                
                r_data[22454] <= r_data[22453];
                
                r_data[22455] <= r_data[22454];
                
                r_data[22456] <= r_data[22455];
                
                r_data[22457] <= r_data[22456];
                
                r_data[22458] <= r_data[22457];
                
                r_data[22459] <= r_data[22458];
                
                r_data[22460] <= r_data[22459];
                
                r_data[22461] <= r_data[22460];
                
                r_data[22462] <= r_data[22461];
                
                r_data[22463] <= r_data[22462];
                
                r_data[22464] <= r_data[22463];
                
                r_data[22465] <= r_data[22464];
                
                r_data[22466] <= r_data[22465];
                
                r_data[22467] <= r_data[22466];
                
                r_data[22468] <= r_data[22467];
                
                r_data[22469] <= r_data[22468];
                
                r_data[22470] <= r_data[22469];
                
                r_data[22471] <= r_data[22470];
                
                r_data[22472] <= r_data[22471];
                
                r_data[22473] <= r_data[22472];
                
                r_data[22474] <= r_data[22473];
                
                r_data[22475] <= r_data[22474];
                
                r_data[22476] <= r_data[22475];
                
                r_data[22477] <= r_data[22476];
                
                r_data[22478] <= r_data[22477];
                
                r_data[22479] <= r_data[22478];
                
                r_data[22480] <= r_data[22479];
                
                r_data[22481] <= r_data[22480];
                
                r_data[22482] <= r_data[22481];
                
                r_data[22483] <= r_data[22482];
                
                r_data[22484] <= r_data[22483];
                
                r_data[22485] <= r_data[22484];
                
                r_data[22486] <= r_data[22485];
                
                r_data[22487] <= r_data[22486];
                
                r_data[22488] <= r_data[22487];
                
                r_data[22489] <= r_data[22488];
                
                r_data[22490] <= r_data[22489];
                
                r_data[22491] <= r_data[22490];
                
                r_data[22492] <= r_data[22491];
                
                r_data[22493] <= r_data[22492];
                
                r_data[22494] <= r_data[22493];
                
                r_data[22495] <= r_data[22494];
                
                r_data[22496] <= r_data[22495];
                
                r_data[22497] <= r_data[22496];
                
                r_data[22498] <= r_data[22497];
                
                r_data[22499] <= r_data[22498];
                
                r_data[22500] <= r_data[22499];
                
                r_data[22501] <= r_data[22500];
                
                r_data[22502] <= r_data[22501];
                
                r_data[22503] <= r_data[22502];
                
                r_data[22504] <= r_data[22503];
                
                r_data[22505] <= r_data[22504];
                
                r_data[22506] <= r_data[22505];
                
                r_data[22507] <= r_data[22506];
                
                r_data[22508] <= r_data[22507];
                
                r_data[22509] <= r_data[22508];
                
                r_data[22510] <= r_data[22509];
                
                r_data[22511] <= r_data[22510];
                
                r_data[22512] <= r_data[22511];
                
                r_data[22513] <= r_data[22512];
                
                r_data[22514] <= r_data[22513];
                
                r_data[22515] <= r_data[22514];
                
                r_data[22516] <= r_data[22515];
                
                r_data[22517] <= r_data[22516];
                
                r_data[22518] <= r_data[22517];
                
                r_data[22519] <= r_data[22518];
                
                r_data[22520] <= r_data[22519];
                
                r_data[22521] <= r_data[22520];
                
                r_data[22522] <= r_data[22521];
                
                r_data[22523] <= r_data[22522];
                
                r_data[22524] <= r_data[22523];
                
                r_data[22525] <= r_data[22524];
                
                r_data[22526] <= r_data[22525];
                
                r_data[22527] <= r_data[22526];
                
                r_data[22528] <= r_data[22527];
                
                r_data[22529] <= r_data[22528];
                
                r_data[22530] <= r_data[22529];
                
                r_data[22531] <= r_data[22530];
                
                r_data[22532] <= r_data[22531];
                
                r_data[22533] <= r_data[22532];
                
                r_data[22534] <= r_data[22533];
                
                r_data[22535] <= r_data[22534];
                
                r_data[22536] <= r_data[22535];
                
                r_data[22537] <= r_data[22536];
                
                r_data[22538] <= r_data[22537];
                
                r_data[22539] <= r_data[22538];
                
                r_data[22540] <= r_data[22539];
                
                r_data[22541] <= r_data[22540];
                
                r_data[22542] <= r_data[22541];
                
                r_data[22543] <= r_data[22542];
                
                r_data[22544] <= r_data[22543];
                
                r_data[22545] <= r_data[22544];
                
                r_data[22546] <= r_data[22545];
                
                r_data[22547] <= r_data[22546];
                
                r_data[22548] <= r_data[22547];
                
                r_data[22549] <= r_data[22548];
                
                r_data[22550] <= r_data[22549];
                
                r_data[22551] <= r_data[22550];
                
                r_data[22552] <= r_data[22551];
                
                r_data[22553] <= r_data[22552];
                
                r_data[22554] <= r_data[22553];
                
                r_data[22555] <= r_data[22554];
                
                r_data[22556] <= r_data[22555];
                
                r_data[22557] <= r_data[22556];
                
                r_data[22558] <= r_data[22557];
                
                r_data[22559] <= r_data[22558];
                
                r_data[22560] <= r_data[22559];
                
                r_data[22561] <= r_data[22560];
                
                r_data[22562] <= r_data[22561];
                
                r_data[22563] <= r_data[22562];
                
                r_data[22564] <= r_data[22563];
                
                r_data[22565] <= r_data[22564];
                
                r_data[22566] <= r_data[22565];
                
                r_data[22567] <= r_data[22566];
                
                r_data[22568] <= r_data[22567];
                
                r_data[22569] <= r_data[22568];
                
                r_data[22570] <= r_data[22569];
                
                r_data[22571] <= r_data[22570];
                
                r_data[22572] <= r_data[22571];
                
                r_data[22573] <= r_data[22572];
                
                r_data[22574] <= r_data[22573];
                
                r_data[22575] <= r_data[22574];
                
                r_data[22576] <= r_data[22575];
                
                r_data[22577] <= r_data[22576];
                
                r_data[22578] <= r_data[22577];
                
                r_data[22579] <= r_data[22578];
                
                r_data[22580] <= r_data[22579];
                
                r_data[22581] <= r_data[22580];
                
                r_data[22582] <= r_data[22581];
                
                r_data[22583] <= r_data[22582];
                
                r_data[22584] <= r_data[22583];
                
                r_data[22585] <= r_data[22584];
                
                r_data[22586] <= r_data[22585];
                
                r_data[22587] <= r_data[22586];
                
                r_data[22588] <= r_data[22587];
                
                r_data[22589] <= r_data[22588];
                
                r_data[22590] <= r_data[22589];
                
                r_data[22591] <= r_data[22590];
                
                r_data[22592] <= r_data[22591];
                
                r_data[22593] <= r_data[22592];
                
                r_data[22594] <= r_data[22593];
                
                r_data[22595] <= r_data[22594];
                
                r_data[22596] <= r_data[22595];
                
                r_data[22597] <= r_data[22596];
                
                r_data[22598] <= r_data[22597];
                
                r_data[22599] <= r_data[22598];
                
                r_data[22600] <= r_data[22599];
                
                r_data[22601] <= r_data[22600];
                
                r_data[22602] <= r_data[22601];
                
                r_data[22603] <= r_data[22602];
                
                r_data[22604] <= r_data[22603];
                
                r_data[22605] <= r_data[22604];
                
                r_data[22606] <= r_data[22605];
                
                r_data[22607] <= r_data[22606];
                
                r_data[22608] <= r_data[22607];
                
                r_data[22609] <= r_data[22608];
                
                r_data[22610] <= r_data[22609];
                
                r_data[22611] <= r_data[22610];
                
                r_data[22612] <= r_data[22611];
                
                r_data[22613] <= r_data[22612];
                
                r_data[22614] <= r_data[22613];
                
                r_data[22615] <= r_data[22614];
                
                r_data[22616] <= r_data[22615];
                
                r_data[22617] <= r_data[22616];
                
                r_data[22618] <= r_data[22617];
                
                r_data[22619] <= r_data[22618];
                
                r_data[22620] <= r_data[22619];
                
                r_data[22621] <= r_data[22620];
                
                r_data[22622] <= r_data[22621];
                
                r_data[22623] <= r_data[22622];
                
                r_data[22624] <= r_data[22623];
                
                r_data[22625] <= r_data[22624];
                
                r_data[22626] <= r_data[22625];
                
                r_data[22627] <= r_data[22626];
                
                r_data[22628] <= r_data[22627];
                
                r_data[22629] <= r_data[22628];
                
                r_data[22630] <= r_data[22629];
                
                r_data[22631] <= r_data[22630];
                
                r_data[22632] <= r_data[22631];
                
                r_data[22633] <= r_data[22632];
                
                r_data[22634] <= r_data[22633];
                
                r_data[22635] <= r_data[22634];
                
                r_data[22636] <= r_data[22635];
                
                r_data[22637] <= r_data[22636];
                
                r_data[22638] <= r_data[22637];
                
                r_data[22639] <= r_data[22638];
                
                r_data[22640] <= r_data[22639];
                
                r_data[22641] <= r_data[22640];
                
                r_data[22642] <= r_data[22641];
                
                r_data[22643] <= r_data[22642];
                
                r_data[22644] <= r_data[22643];
                
                r_data[22645] <= r_data[22644];
                
                r_data[22646] <= r_data[22645];
                
                r_data[22647] <= r_data[22646];
                
                r_data[22648] <= r_data[22647];
                
                r_data[22649] <= r_data[22648];
                
                r_data[22650] <= r_data[22649];
                
                r_data[22651] <= r_data[22650];
                
                r_data[22652] <= r_data[22651];
                
                r_data[22653] <= r_data[22652];
                
                r_data[22654] <= r_data[22653];
                
                r_data[22655] <= r_data[22654];
                
                r_data[22656] <= r_data[22655];
                
                r_data[22657] <= r_data[22656];
                
                r_data[22658] <= r_data[22657];
                
                r_data[22659] <= r_data[22658];
                
                r_data[22660] <= r_data[22659];
                
                r_data[22661] <= r_data[22660];
                
                r_data[22662] <= r_data[22661];
                
                r_data[22663] <= r_data[22662];
                
                r_data[22664] <= r_data[22663];
                
                r_data[22665] <= r_data[22664];
                
                r_data[22666] <= r_data[22665];
                
                r_data[22667] <= r_data[22666];
                
                r_data[22668] <= r_data[22667];
                
                r_data[22669] <= r_data[22668];
                
                r_data[22670] <= r_data[22669];
                
                r_data[22671] <= r_data[22670];
                
                r_data[22672] <= r_data[22671];
                
                r_data[22673] <= r_data[22672];
                
                r_data[22674] <= r_data[22673];
                
                r_data[22675] <= r_data[22674];
                
                r_data[22676] <= r_data[22675];
                
                r_data[22677] <= r_data[22676];
                
                r_data[22678] <= r_data[22677];
                
                r_data[22679] <= r_data[22678];
                
                r_data[22680] <= r_data[22679];
                
                r_data[22681] <= r_data[22680];
                
                r_data[22682] <= r_data[22681];
                
                r_data[22683] <= r_data[22682];
                
                r_data[22684] <= r_data[22683];
                
                r_data[22685] <= r_data[22684];
                
                r_data[22686] <= r_data[22685];
                
                r_data[22687] <= r_data[22686];
                
                r_data[22688] <= r_data[22687];
                
                r_data[22689] <= r_data[22688];
                
                r_data[22690] <= r_data[22689];
                
                r_data[22691] <= r_data[22690];
                
                r_data[22692] <= r_data[22691];
                
                r_data[22693] <= r_data[22692];
                
                r_data[22694] <= r_data[22693];
                
                r_data[22695] <= r_data[22694];
                
                r_data[22696] <= r_data[22695];
                
                r_data[22697] <= r_data[22696];
                
                r_data[22698] <= r_data[22697];
                
                r_data[22699] <= r_data[22698];
                
                r_data[22700] <= r_data[22699];
                
                r_data[22701] <= r_data[22700];
                
                r_data[22702] <= r_data[22701];
                
                r_data[22703] <= r_data[22702];
                
                r_data[22704] <= r_data[22703];
                
                r_data[22705] <= r_data[22704];
                
                r_data[22706] <= r_data[22705];
                
                r_data[22707] <= r_data[22706];
                
                r_data[22708] <= r_data[22707];
                
                r_data[22709] <= r_data[22708];
                
                r_data[22710] <= r_data[22709];
                
                r_data[22711] <= r_data[22710];
                
                r_data[22712] <= r_data[22711];
                
                r_data[22713] <= r_data[22712];
                
                r_data[22714] <= r_data[22713];
                
                r_data[22715] <= r_data[22714];
                
                r_data[22716] <= r_data[22715];
                
                r_data[22717] <= r_data[22716];
                
                r_data[22718] <= r_data[22717];
                
                r_data[22719] <= r_data[22718];
                
                r_data[22720] <= r_data[22719];
                
                r_data[22721] <= r_data[22720];
                
                r_data[22722] <= r_data[22721];
                
                r_data[22723] <= r_data[22722];
                
                r_data[22724] <= r_data[22723];
                
                r_data[22725] <= r_data[22724];
                
                r_data[22726] <= r_data[22725];
                
                r_data[22727] <= r_data[22726];
                
                r_data[22728] <= r_data[22727];
                
                r_data[22729] <= r_data[22728];
                
                r_data[22730] <= r_data[22729];
                
                r_data[22731] <= r_data[22730];
                
                r_data[22732] <= r_data[22731];
                
                r_data[22733] <= r_data[22732];
                
                r_data[22734] <= r_data[22733];
                
                r_data[22735] <= r_data[22734];
                
                r_data[22736] <= r_data[22735];
                
                r_data[22737] <= r_data[22736];
                
                r_data[22738] <= r_data[22737];
                
                r_data[22739] <= r_data[22738];
                
                r_data[22740] <= r_data[22739];
                
                r_data[22741] <= r_data[22740];
                
                r_data[22742] <= r_data[22741];
                
                r_data[22743] <= r_data[22742];
                
                r_data[22744] <= r_data[22743];
                
                r_data[22745] <= r_data[22744];
                
                r_data[22746] <= r_data[22745];
                
                r_data[22747] <= r_data[22746];
                
                r_data[22748] <= r_data[22747];
                
                r_data[22749] <= r_data[22748];
                
                r_data[22750] <= r_data[22749];
                
                r_data[22751] <= r_data[22750];
                
                r_data[22752] <= r_data[22751];
                
                r_data[22753] <= r_data[22752];
                
                r_data[22754] <= r_data[22753];
                
                r_data[22755] <= r_data[22754];
                
                r_data[22756] <= r_data[22755];
                
                r_data[22757] <= r_data[22756];
                
                r_data[22758] <= r_data[22757];
                
                r_data[22759] <= r_data[22758];
                
                r_data[22760] <= r_data[22759];
                
                r_data[22761] <= r_data[22760];
                
                r_data[22762] <= r_data[22761];
                
                r_data[22763] <= r_data[22762];
                
                r_data[22764] <= r_data[22763];
                
                r_data[22765] <= r_data[22764];
                
                r_data[22766] <= r_data[22765];
                
                r_data[22767] <= r_data[22766];
                
                r_data[22768] <= r_data[22767];
                
                r_data[22769] <= r_data[22768];
                
                r_data[22770] <= r_data[22769];
                
                r_data[22771] <= r_data[22770];
                
                r_data[22772] <= r_data[22771];
                
                r_data[22773] <= r_data[22772];
                
                r_data[22774] <= r_data[22773];
                
                r_data[22775] <= r_data[22774];
                
                r_data[22776] <= r_data[22775];
                
                r_data[22777] <= r_data[22776];
                
                r_data[22778] <= r_data[22777];
                
                r_data[22779] <= r_data[22778];
                
                r_data[22780] <= r_data[22779];
                
                r_data[22781] <= r_data[22780];
                
                r_data[22782] <= r_data[22781];
                
                r_data[22783] <= r_data[22782];
                
                r_data[22784] <= r_data[22783];
                
                r_data[22785] <= r_data[22784];
                
                r_data[22786] <= r_data[22785];
                
                r_data[22787] <= r_data[22786];
                
                r_data[22788] <= r_data[22787];
                
                r_data[22789] <= r_data[22788];
                
                r_data[22790] <= r_data[22789];
                
                r_data[22791] <= r_data[22790];
                
                r_data[22792] <= r_data[22791];
                
                r_data[22793] <= r_data[22792];
                
                r_data[22794] <= r_data[22793];
                
                r_data[22795] <= r_data[22794];
                
                r_data[22796] <= r_data[22795];
                
                r_data[22797] <= r_data[22796];
                
                r_data[22798] <= r_data[22797];
                
                r_data[22799] <= r_data[22798];
                
                r_data[22800] <= r_data[22799];
                
                r_data[22801] <= r_data[22800];
                
                r_data[22802] <= r_data[22801];
                
                r_data[22803] <= r_data[22802];
                
                r_data[22804] <= r_data[22803];
                
                r_data[22805] <= r_data[22804];
                
                r_data[22806] <= r_data[22805];
                
                r_data[22807] <= r_data[22806];
                
                r_data[22808] <= r_data[22807];
                
                r_data[22809] <= r_data[22808];
                
                r_data[22810] <= r_data[22809];
                
                r_data[22811] <= r_data[22810];
                
                r_data[22812] <= r_data[22811];
                
                r_data[22813] <= r_data[22812];
                
                r_data[22814] <= r_data[22813];
                
                r_data[22815] <= r_data[22814];
                
                r_data[22816] <= r_data[22815];
                
                r_data[22817] <= r_data[22816];
                
                r_data[22818] <= r_data[22817];
                
                r_data[22819] <= r_data[22818];
                
                r_data[22820] <= r_data[22819];
                
                r_data[22821] <= r_data[22820];
                
                r_data[22822] <= r_data[22821];
                
                r_data[22823] <= r_data[22822];
                
                r_data[22824] <= r_data[22823];
                
                r_data[22825] <= r_data[22824];
                
                r_data[22826] <= r_data[22825];
                
                r_data[22827] <= r_data[22826];
                
                r_data[22828] <= r_data[22827];
                
                r_data[22829] <= r_data[22828];
                
                r_data[22830] <= r_data[22829];
                
                r_data[22831] <= r_data[22830];
                
                r_data[22832] <= r_data[22831];
                
                r_data[22833] <= r_data[22832];
                
                r_data[22834] <= r_data[22833];
                
                r_data[22835] <= r_data[22834];
                
                r_data[22836] <= r_data[22835];
                
                r_data[22837] <= r_data[22836];
                
                r_data[22838] <= r_data[22837];
                
                r_data[22839] <= r_data[22838];
                
                r_data[22840] <= r_data[22839];
                
                r_data[22841] <= r_data[22840];
                
                r_data[22842] <= r_data[22841];
                
                r_data[22843] <= r_data[22842];
                
                r_data[22844] <= r_data[22843];
                
                r_data[22845] <= r_data[22844];
                
                r_data[22846] <= r_data[22845];
                
                r_data[22847] <= r_data[22846];
                
                r_data[22848] <= r_data[22847];
                
                r_data[22849] <= r_data[22848];
                
                r_data[22850] <= r_data[22849];
                
                r_data[22851] <= r_data[22850];
                
                r_data[22852] <= r_data[22851];
                
                r_data[22853] <= r_data[22852];
                
                r_data[22854] <= r_data[22853];
                
                r_data[22855] <= r_data[22854];
                
                r_data[22856] <= r_data[22855];
                
                r_data[22857] <= r_data[22856];
                
                r_data[22858] <= r_data[22857];
                
                r_data[22859] <= r_data[22858];
                
                r_data[22860] <= r_data[22859];
                
                r_data[22861] <= r_data[22860];
                
                r_data[22862] <= r_data[22861];
                
                r_data[22863] <= r_data[22862];
                
                r_data[22864] <= r_data[22863];
                
                r_data[22865] <= r_data[22864];
                
                r_data[22866] <= r_data[22865];
                
                r_data[22867] <= r_data[22866];
                
                r_data[22868] <= r_data[22867];
                
                r_data[22869] <= r_data[22868];
                
                r_data[22870] <= r_data[22869];
                
                r_data[22871] <= r_data[22870];
                
                r_data[22872] <= r_data[22871];
                
                r_data[22873] <= r_data[22872];
                
                r_data[22874] <= r_data[22873];
                
                r_data[22875] <= r_data[22874];
                
                r_data[22876] <= r_data[22875];
                
                r_data[22877] <= r_data[22876];
                
                r_data[22878] <= r_data[22877];
                
                r_data[22879] <= r_data[22878];
                
                r_data[22880] <= r_data[22879];
                
                r_data[22881] <= r_data[22880];
                
                r_data[22882] <= r_data[22881];
                
                r_data[22883] <= r_data[22882];
                
                r_data[22884] <= r_data[22883];
                
                r_data[22885] <= r_data[22884];
                
                r_data[22886] <= r_data[22885];
                
                r_data[22887] <= r_data[22886];
                
                r_data[22888] <= r_data[22887];
                
                r_data[22889] <= r_data[22888];
                
                r_data[22890] <= r_data[22889];
                
                r_data[22891] <= r_data[22890];
                
                r_data[22892] <= r_data[22891];
                
                r_data[22893] <= r_data[22892];
                
                r_data[22894] <= r_data[22893];
                
                r_data[22895] <= r_data[22894];
                
                r_data[22896] <= r_data[22895];
                
                r_data[22897] <= r_data[22896];
                
                r_data[22898] <= r_data[22897];
                
                r_data[22899] <= r_data[22898];
                
                r_data[22900] <= r_data[22899];
                
                r_data[22901] <= r_data[22900];
                
                r_data[22902] <= r_data[22901];
                
                r_data[22903] <= r_data[22902];
                
                r_data[22904] <= r_data[22903];
                
                r_data[22905] <= r_data[22904];
                
                r_data[22906] <= r_data[22905];
                
                r_data[22907] <= r_data[22906];
                
                r_data[22908] <= r_data[22907];
                
                r_data[22909] <= r_data[22908];
                
                r_data[22910] <= r_data[22909];
                
                r_data[22911] <= r_data[22910];
                
                r_data[22912] <= r_data[22911];
                
                r_data[22913] <= r_data[22912];
                
                r_data[22914] <= r_data[22913];
                
                r_data[22915] <= r_data[22914];
                
                r_data[22916] <= r_data[22915];
                
                r_data[22917] <= r_data[22916];
                
                r_data[22918] <= r_data[22917];
                
                r_data[22919] <= r_data[22918];
                
                r_data[22920] <= r_data[22919];
                
                r_data[22921] <= r_data[22920];
                
                r_data[22922] <= r_data[22921];
                
                r_data[22923] <= r_data[22922];
                
                r_data[22924] <= r_data[22923];
                
                r_data[22925] <= r_data[22924];
                
                r_data[22926] <= r_data[22925];
                
                r_data[22927] <= r_data[22926];
                
                r_data[22928] <= r_data[22927];
                
                r_data[22929] <= r_data[22928];
                
                r_data[22930] <= r_data[22929];
                
                r_data[22931] <= r_data[22930];
                
                r_data[22932] <= r_data[22931];
                
                r_data[22933] <= r_data[22932];
                
                r_data[22934] <= r_data[22933];
                
                r_data[22935] <= r_data[22934];
                
                r_data[22936] <= r_data[22935];
                
                r_data[22937] <= r_data[22936];
                
                r_data[22938] <= r_data[22937];
                
                r_data[22939] <= r_data[22938];
                
                r_data[22940] <= r_data[22939];
                
                r_data[22941] <= r_data[22940];
                
                r_data[22942] <= r_data[22941];
                
                r_data[22943] <= r_data[22942];
                
                r_data[22944] <= r_data[22943];
                
                r_data[22945] <= r_data[22944];
                
                r_data[22946] <= r_data[22945];
                
                r_data[22947] <= r_data[22946];
                
                r_data[22948] <= r_data[22947];
                
                r_data[22949] <= r_data[22948];
                
                r_data[22950] <= r_data[22949];
                
                r_data[22951] <= r_data[22950];
                
                r_data[22952] <= r_data[22951];
                
                r_data[22953] <= r_data[22952];
                
                r_data[22954] <= r_data[22953];
                
                r_data[22955] <= r_data[22954];
                
                r_data[22956] <= r_data[22955];
                
                r_data[22957] <= r_data[22956];
                
                r_data[22958] <= r_data[22957];
                
                r_data[22959] <= r_data[22958];
                
                r_data[22960] <= r_data[22959];
                
                r_data[22961] <= r_data[22960];
                
                r_data[22962] <= r_data[22961];
                
                r_data[22963] <= r_data[22962];
                
                r_data[22964] <= r_data[22963];
                
                r_data[22965] <= r_data[22964];
                
                r_data[22966] <= r_data[22965];
                
                r_data[22967] <= r_data[22966];
                
                r_data[22968] <= r_data[22967];
                
                r_data[22969] <= r_data[22968];
                
                r_data[22970] <= r_data[22969];
                
                r_data[22971] <= r_data[22970];
                
                r_data[22972] <= r_data[22971];
                
                r_data[22973] <= r_data[22972];
                
                r_data[22974] <= r_data[22973];
                
                r_data[22975] <= r_data[22974];
                
                r_data[22976] <= r_data[22975];
                
                r_data[22977] <= r_data[22976];
                
                r_data[22978] <= r_data[22977];
                
                r_data[22979] <= r_data[22978];
                
                r_data[22980] <= r_data[22979];
                
                r_data[22981] <= r_data[22980];
                
                r_data[22982] <= r_data[22981];
                
                r_data[22983] <= r_data[22982];
                
                r_data[22984] <= r_data[22983];
                
                r_data[22985] <= r_data[22984];
                
                r_data[22986] <= r_data[22985];
                
                r_data[22987] <= r_data[22986];
                
                r_data[22988] <= r_data[22987];
                
                r_data[22989] <= r_data[22988];
                
                r_data[22990] <= r_data[22989];
                
                r_data[22991] <= r_data[22990];
                
                r_data[22992] <= r_data[22991];
                
                r_data[22993] <= r_data[22992];
                
                r_data[22994] <= r_data[22993];
                
                r_data[22995] <= r_data[22994];
                
                r_data[22996] <= r_data[22995];
                
                r_data[22997] <= r_data[22996];
                
                r_data[22998] <= r_data[22997];
                
                r_data[22999] <= r_data[22998];
                
                r_data[23000] <= r_data[22999];
                
                r_data[23001] <= r_data[23000];
                
                r_data[23002] <= r_data[23001];
                
                r_data[23003] <= r_data[23002];
                
                r_data[23004] <= r_data[23003];
                
                r_data[23005] <= r_data[23004];
                
                r_data[23006] <= r_data[23005];
                
                r_data[23007] <= r_data[23006];
                
                r_data[23008] <= r_data[23007];
                
                r_data[23009] <= r_data[23008];
                
                r_data[23010] <= r_data[23009];
                
                r_data[23011] <= r_data[23010];
                
                r_data[23012] <= r_data[23011];
                
                r_data[23013] <= r_data[23012];
                
                r_data[23014] <= r_data[23013];
                
                r_data[23015] <= r_data[23014];
                
                r_data[23016] <= r_data[23015];
                
                r_data[23017] <= r_data[23016];
                
                r_data[23018] <= r_data[23017];
                
                r_data[23019] <= r_data[23018];
                
                r_data[23020] <= r_data[23019];
                
                r_data[23021] <= r_data[23020];
                
                r_data[23022] <= r_data[23021];
                
                r_data[23023] <= r_data[23022];
                
                r_data[23024] <= r_data[23023];
                
                r_data[23025] <= r_data[23024];
                
                r_data[23026] <= r_data[23025];
                
                r_data[23027] <= r_data[23026];
                
                r_data[23028] <= r_data[23027];
                
                r_data[23029] <= r_data[23028];
                
                r_data[23030] <= r_data[23029];
                
                r_data[23031] <= r_data[23030];
                
                r_data[23032] <= r_data[23031];
                
                r_data[23033] <= r_data[23032];
                
                r_data[23034] <= r_data[23033];
                
                r_data[23035] <= r_data[23034];
                
                r_data[23036] <= r_data[23035];
                
                r_data[23037] <= r_data[23036];
                
                r_data[23038] <= r_data[23037];
                
                r_data[23039] <= r_data[23038];
                
                r_data[23040] <= r_data[23039];
                
                r_data[23041] <= r_data[23040];
                
                r_data[23042] <= r_data[23041];
                
                r_data[23043] <= r_data[23042];
                
                r_data[23044] <= r_data[23043];
                
                r_data[23045] <= r_data[23044];
                
                r_data[23046] <= r_data[23045];
                
                r_data[23047] <= r_data[23046];
                
                r_data[23048] <= r_data[23047];
                
                r_data[23049] <= r_data[23048];
                
                r_data[23050] <= r_data[23049];
                
                r_data[23051] <= r_data[23050];
                
                r_data[23052] <= r_data[23051];
                
                r_data[23053] <= r_data[23052];
                
                r_data[23054] <= r_data[23053];
                
                r_data[23055] <= r_data[23054];
                
                r_data[23056] <= r_data[23055];
                
                r_data[23057] <= r_data[23056];
                
                r_data[23058] <= r_data[23057];
                
                r_data[23059] <= r_data[23058];
                
                r_data[23060] <= r_data[23059];
                
                r_data[23061] <= r_data[23060];
                
                r_data[23062] <= r_data[23061];
                
                r_data[23063] <= r_data[23062];
                
                r_data[23064] <= r_data[23063];
                
                r_data[23065] <= r_data[23064];
                
                r_data[23066] <= r_data[23065];
                
                r_data[23067] <= r_data[23066];
                
                r_data[23068] <= r_data[23067];
                
                r_data[23069] <= r_data[23068];
                
                r_data[23070] <= r_data[23069];
                
                r_data[23071] <= r_data[23070];
                
                r_data[23072] <= r_data[23071];
                
                r_data[23073] <= r_data[23072];
                
                r_data[23074] <= r_data[23073];
                
                r_data[23075] <= r_data[23074];
                
                r_data[23076] <= r_data[23075];
                
                r_data[23077] <= r_data[23076];
                
                r_data[23078] <= r_data[23077];
                
                r_data[23079] <= r_data[23078];
                
                r_data[23080] <= r_data[23079];
                
                r_data[23081] <= r_data[23080];
                
                r_data[23082] <= r_data[23081];
                
                r_data[23083] <= r_data[23082];
                
                r_data[23084] <= r_data[23083];
                
                r_data[23085] <= r_data[23084];
                
                r_data[23086] <= r_data[23085];
                
                r_data[23087] <= r_data[23086];
                
                r_data[23088] <= r_data[23087];
                
                r_data[23089] <= r_data[23088];
                
                r_data[23090] <= r_data[23089];
                
                r_data[23091] <= r_data[23090];
                
                r_data[23092] <= r_data[23091];
                
                r_data[23093] <= r_data[23092];
                
                r_data[23094] <= r_data[23093];
                
                r_data[23095] <= r_data[23094];
                
                r_data[23096] <= r_data[23095];
                
                r_data[23097] <= r_data[23096];
                
                r_data[23098] <= r_data[23097];
                
                r_data[23099] <= r_data[23098];
                
                r_data[23100] <= r_data[23099];
                
                r_data[23101] <= r_data[23100];
                
                r_data[23102] <= r_data[23101];
                
                r_data[23103] <= r_data[23102];
                
                r_data[23104] <= r_data[23103];
                
                r_data[23105] <= r_data[23104];
                
                r_data[23106] <= r_data[23105];
                
                r_data[23107] <= r_data[23106];
                
                r_data[23108] <= r_data[23107];
                
                r_data[23109] <= r_data[23108];
                
                r_data[23110] <= r_data[23109];
                
                r_data[23111] <= r_data[23110];
                
                r_data[23112] <= r_data[23111];
                
                r_data[23113] <= r_data[23112];
                
                r_data[23114] <= r_data[23113];
                
                r_data[23115] <= r_data[23114];
                
                r_data[23116] <= r_data[23115];
                
                r_data[23117] <= r_data[23116];
                
                r_data[23118] <= r_data[23117];
                
                r_data[23119] <= r_data[23118];
                
                r_data[23120] <= r_data[23119];
                
                r_data[23121] <= r_data[23120];
                
                r_data[23122] <= r_data[23121];
                
                r_data[23123] <= r_data[23122];
                
                r_data[23124] <= r_data[23123];
                
                r_data[23125] <= r_data[23124];
                
                r_data[23126] <= r_data[23125];
                
                r_data[23127] <= r_data[23126];
                
                r_data[23128] <= r_data[23127];
                
                r_data[23129] <= r_data[23128];
                
                r_data[23130] <= r_data[23129];
                
                r_data[23131] <= r_data[23130];
                
                r_data[23132] <= r_data[23131];
                
                r_data[23133] <= r_data[23132];
                
                r_data[23134] <= r_data[23133];
                
                r_data[23135] <= r_data[23134];
                
                r_data[23136] <= r_data[23135];
                
                r_data[23137] <= r_data[23136];
                
                r_data[23138] <= r_data[23137];
                
                r_data[23139] <= r_data[23138];
                
                r_data[23140] <= r_data[23139];
                
                r_data[23141] <= r_data[23140];
                
                r_data[23142] <= r_data[23141];
                
                r_data[23143] <= r_data[23142];
                
                r_data[23144] <= r_data[23143];
                
                r_data[23145] <= r_data[23144];
                
                r_data[23146] <= r_data[23145];
                
                r_data[23147] <= r_data[23146];
                
                r_data[23148] <= r_data[23147];
                
                r_data[23149] <= r_data[23148];
                
                r_data[23150] <= r_data[23149];
                
                r_data[23151] <= r_data[23150];
                
                r_data[23152] <= r_data[23151];
                
                r_data[23153] <= r_data[23152];
                
                r_data[23154] <= r_data[23153];
                
                r_data[23155] <= r_data[23154];
                
                r_data[23156] <= r_data[23155];
                
                r_data[23157] <= r_data[23156];
                
                r_data[23158] <= r_data[23157];
                
                r_data[23159] <= r_data[23158];
                
                r_data[23160] <= r_data[23159];
                
                r_data[23161] <= r_data[23160];
                
                r_data[23162] <= r_data[23161];
                
                r_data[23163] <= r_data[23162];
                
                r_data[23164] <= r_data[23163];
                
                r_data[23165] <= r_data[23164];
                
                r_data[23166] <= r_data[23165];
                
                r_data[23167] <= r_data[23166];
                
                r_data[23168] <= r_data[23167];
                
                r_data[23169] <= r_data[23168];
                
                r_data[23170] <= r_data[23169];
                
                r_data[23171] <= r_data[23170];
                
                r_data[23172] <= r_data[23171];
                
                r_data[23173] <= r_data[23172];
                
                r_data[23174] <= r_data[23173];
                
                r_data[23175] <= r_data[23174];
                
                r_data[23176] <= r_data[23175];
                
                r_data[23177] <= r_data[23176];
                
                r_data[23178] <= r_data[23177];
                
                r_data[23179] <= r_data[23178];
                
                r_data[23180] <= r_data[23179];
                
                r_data[23181] <= r_data[23180];
                
                r_data[23182] <= r_data[23181];
                
                r_data[23183] <= r_data[23182];
                
                r_data[23184] <= r_data[23183];
                
                r_data[23185] <= r_data[23184];
                
                r_data[23186] <= r_data[23185];
                
                r_data[23187] <= r_data[23186];
                
                r_data[23188] <= r_data[23187];
                
                r_data[23189] <= r_data[23188];
                
                r_data[23190] <= r_data[23189];
                
                r_data[23191] <= r_data[23190];
                
                r_data[23192] <= r_data[23191];
                
                r_data[23193] <= r_data[23192];
                
                r_data[23194] <= r_data[23193];
                
                r_data[23195] <= r_data[23194];
                
                r_data[23196] <= r_data[23195];
                
                r_data[23197] <= r_data[23196];
                
                r_data[23198] <= r_data[23197];
                
                r_data[23199] <= r_data[23198];
                
                r_data[23200] <= r_data[23199];
                
                r_data[23201] <= r_data[23200];
                
                r_data[23202] <= r_data[23201];
                
                r_data[23203] <= r_data[23202];
                
                r_data[23204] <= r_data[23203];
                
                r_data[23205] <= r_data[23204];
                
                r_data[23206] <= r_data[23205];
                
                r_data[23207] <= r_data[23206];
                
                r_data[23208] <= r_data[23207];
                
                r_data[23209] <= r_data[23208];
                
                r_data[23210] <= r_data[23209];
                
                r_data[23211] <= r_data[23210];
                
                r_data[23212] <= r_data[23211];
                
                r_data[23213] <= r_data[23212];
                
                r_data[23214] <= r_data[23213];
                
                r_data[23215] <= r_data[23214];
                
                r_data[23216] <= r_data[23215];
                
                r_data[23217] <= r_data[23216];
                
                r_data[23218] <= r_data[23217];
                
                r_data[23219] <= r_data[23218];
                
                r_data[23220] <= r_data[23219];
                
                r_data[23221] <= r_data[23220];
                
                r_data[23222] <= r_data[23221];
                
                r_data[23223] <= r_data[23222];
                
                r_data[23224] <= r_data[23223];
                
                r_data[23225] <= r_data[23224];
                
                r_data[23226] <= r_data[23225];
                
                r_data[23227] <= r_data[23226];
                
                r_data[23228] <= r_data[23227];
                
                r_data[23229] <= r_data[23228];
                
                r_data[23230] <= r_data[23229];
                
                r_data[23231] <= r_data[23230];
                
                r_data[23232] <= r_data[23231];
                
                r_data[23233] <= r_data[23232];
                
                r_data[23234] <= r_data[23233];
                
                r_data[23235] <= r_data[23234];
                
                r_data[23236] <= r_data[23235];
                
                r_data[23237] <= r_data[23236];
                
                r_data[23238] <= r_data[23237];
                
                r_data[23239] <= r_data[23238];
                
                r_data[23240] <= r_data[23239];
                
                r_data[23241] <= r_data[23240];
                
                r_data[23242] <= r_data[23241];
                
                r_data[23243] <= r_data[23242];
                
                r_data[23244] <= r_data[23243];
                
                r_data[23245] <= r_data[23244];
                
                r_data[23246] <= r_data[23245];
                
                r_data[23247] <= r_data[23246];
                
                r_data[23248] <= r_data[23247];
                
                r_data[23249] <= r_data[23248];
                
                r_data[23250] <= r_data[23249];
                
                r_data[23251] <= r_data[23250];
                
                r_data[23252] <= r_data[23251];
                
                r_data[23253] <= r_data[23252];
                
                r_data[23254] <= r_data[23253];
                
                r_data[23255] <= r_data[23254];
                
                r_data[23256] <= r_data[23255];
                
                r_data[23257] <= r_data[23256];
                
                r_data[23258] <= r_data[23257];
                
                r_data[23259] <= r_data[23258];
                
                r_data[23260] <= r_data[23259];
                
                r_data[23261] <= r_data[23260];
                
                r_data[23262] <= r_data[23261];
                
                r_data[23263] <= r_data[23262];
                
                r_data[23264] <= r_data[23263];
                
                r_data[23265] <= r_data[23264];
                
                r_data[23266] <= r_data[23265];
                
                r_data[23267] <= r_data[23266];
                
                r_data[23268] <= r_data[23267];
                
                r_data[23269] <= r_data[23268];
                
                r_data[23270] <= r_data[23269];
                
                r_data[23271] <= r_data[23270];
                
                r_data[23272] <= r_data[23271];
                
                r_data[23273] <= r_data[23272];
                
                r_data[23274] <= r_data[23273];
                
                r_data[23275] <= r_data[23274];
                
                r_data[23276] <= r_data[23275];
                
                r_data[23277] <= r_data[23276];
                
                r_data[23278] <= r_data[23277];
                
                r_data[23279] <= r_data[23278];
                
                r_data[23280] <= r_data[23279];
                
                r_data[23281] <= r_data[23280];
                
                r_data[23282] <= r_data[23281];
                
                r_data[23283] <= r_data[23282];
                
                r_data[23284] <= r_data[23283];
                
                r_data[23285] <= r_data[23284];
                
                r_data[23286] <= r_data[23285];
                
                r_data[23287] <= r_data[23286];
                
                r_data[23288] <= r_data[23287];
                
                r_data[23289] <= r_data[23288];
                
                r_data[23290] <= r_data[23289];
                
                r_data[23291] <= r_data[23290];
                
                r_data[23292] <= r_data[23291];
                
                r_data[23293] <= r_data[23292];
                
                r_data[23294] <= r_data[23293];
                
                r_data[23295] <= r_data[23294];
                
                r_data[23296] <= r_data[23295];
                
                r_data[23297] <= r_data[23296];
                
                r_data[23298] <= r_data[23297];
                
                r_data[23299] <= r_data[23298];
                
                r_data[23300] <= r_data[23299];
                
                r_data[23301] <= r_data[23300];
                
                r_data[23302] <= r_data[23301];
                
                r_data[23303] <= r_data[23302];
                
                r_data[23304] <= r_data[23303];
                
                r_data[23305] <= r_data[23304];
                
                r_data[23306] <= r_data[23305];
                
                r_data[23307] <= r_data[23306];
                
                r_data[23308] <= r_data[23307];
                
                r_data[23309] <= r_data[23308];
                
                r_data[23310] <= r_data[23309];
                
                r_data[23311] <= r_data[23310];
                
                r_data[23312] <= r_data[23311];
                
                r_data[23313] <= r_data[23312];
                
                r_data[23314] <= r_data[23313];
                
                r_data[23315] <= r_data[23314];
                
                r_data[23316] <= r_data[23315];
                
                r_data[23317] <= r_data[23316];
                
                r_data[23318] <= r_data[23317];
                
                r_data[23319] <= r_data[23318];
                
                r_data[23320] <= r_data[23319];
                
                r_data[23321] <= r_data[23320];
                
                r_data[23322] <= r_data[23321];
                
                r_data[23323] <= r_data[23322];
                
                r_data[23324] <= r_data[23323];
                
                r_data[23325] <= r_data[23324];
                
                r_data[23326] <= r_data[23325];
                
                r_data[23327] <= r_data[23326];
                
                r_data[23328] <= r_data[23327];
                
                r_data[23329] <= r_data[23328];
                
                r_data[23330] <= r_data[23329];
                
                r_data[23331] <= r_data[23330];
                
                r_data[23332] <= r_data[23331];
                
                r_data[23333] <= r_data[23332];
                
                r_data[23334] <= r_data[23333];
                
                r_data[23335] <= r_data[23334];
                
                r_data[23336] <= r_data[23335];
                
                r_data[23337] <= r_data[23336];
                
                r_data[23338] <= r_data[23337];
                
                r_data[23339] <= r_data[23338];
                
                r_data[23340] <= r_data[23339];
                
                r_data[23341] <= r_data[23340];
                
                r_data[23342] <= r_data[23341];
                
                r_data[23343] <= r_data[23342];
                
                r_data[23344] <= r_data[23343];
                
                r_data[23345] <= r_data[23344];
                
                r_data[23346] <= r_data[23345];
                
                r_data[23347] <= r_data[23346];
                
                r_data[23348] <= r_data[23347];
                
                r_data[23349] <= r_data[23348];
                
                r_data[23350] <= r_data[23349];
                
                r_data[23351] <= r_data[23350];
                
                r_data[23352] <= r_data[23351];
                
                r_data[23353] <= r_data[23352];
                
                r_data[23354] <= r_data[23353];
                
                r_data[23355] <= r_data[23354];
                
                r_data[23356] <= r_data[23355];
                
                r_data[23357] <= r_data[23356];
                
                r_data[23358] <= r_data[23357];
                
                r_data[23359] <= r_data[23358];
                
                r_data[23360] <= r_data[23359];
                
                r_data[23361] <= r_data[23360];
                
                r_data[23362] <= r_data[23361];
                
                r_data[23363] <= r_data[23362];
                
                r_data[23364] <= r_data[23363];
                
                r_data[23365] <= r_data[23364];
                
                r_data[23366] <= r_data[23365];
                
                r_data[23367] <= r_data[23366];
                
                r_data[23368] <= r_data[23367];
                
                r_data[23369] <= r_data[23368];
                
                r_data[23370] <= r_data[23369];
                
                r_data[23371] <= r_data[23370];
                
                r_data[23372] <= r_data[23371];
                
                r_data[23373] <= r_data[23372];
                
                r_data[23374] <= r_data[23373];
                
                r_data[23375] <= r_data[23374];
                
                r_data[23376] <= r_data[23375];
                
                r_data[23377] <= r_data[23376];
                
                r_data[23378] <= r_data[23377];
                
                r_data[23379] <= r_data[23378];
                
                r_data[23380] <= r_data[23379];
                
                r_data[23381] <= r_data[23380];
                
                r_data[23382] <= r_data[23381];
                
                r_data[23383] <= r_data[23382];
                
                r_data[23384] <= r_data[23383];
                
                r_data[23385] <= r_data[23384];
                
                r_data[23386] <= r_data[23385];
                
                r_data[23387] <= r_data[23386];
                
                r_data[23388] <= r_data[23387];
                
                r_data[23389] <= r_data[23388];
                
                r_data[23390] <= r_data[23389];
                
                r_data[23391] <= r_data[23390];
                
                r_data[23392] <= r_data[23391];
                
                r_data[23393] <= r_data[23392];
                
                r_data[23394] <= r_data[23393];
                
                r_data[23395] <= r_data[23394];
                
                r_data[23396] <= r_data[23395];
                
                r_data[23397] <= r_data[23396];
                
                r_data[23398] <= r_data[23397];
                
                r_data[23399] <= r_data[23398];
                
                r_data[23400] <= r_data[23399];
                
                r_data[23401] <= r_data[23400];
                
                r_data[23402] <= r_data[23401];
                
                r_data[23403] <= r_data[23402];
                
                r_data[23404] <= r_data[23403];
                
                r_data[23405] <= r_data[23404];
                
                r_data[23406] <= r_data[23405];
                
                r_data[23407] <= r_data[23406];
                
                r_data[23408] <= r_data[23407];
                
                r_data[23409] <= r_data[23408];
                
                r_data[23410] <= r_data[23409];
                
                r_data[23411] <= r_data[23410];
                
                r_data[23412] <= r_data[23411];
                
                r_data[23413] <= r_data[23412];
                
                r_data[23414] <= r_data[23413];
                
                r_data[23415] <= r_data[23414];
                
                r_data[23416] <= r_data[23415];
                
                r_data[23417] <= r_data[23416];
                
                r_data[23418] <= r_data[23417];
                
                r_data[23419] <= r_data[23418];
                
                r_data[23420] <= r_data[23419];
                
                r_data[23421] <= r_data[23420];
                
                r_data[23422] <= r_data[23421];
                
                r_data[23423] <= r_data[23422];
                
                r_data[23424] <= r_data[23423];
                
                r_data[23425] <= r_data[23424];
                
                r_data[23426] <= r_data[23425];
                
                r_data[23427] <= r_data[23426];
                
                r_data[23428] <= r_data[23427];
                
                r_data[23429] <= r_data[23428];
                
                r_data[23430] <= r_data[23429];
                
                r_data[23431] <= r_data[23430];
                
                r_data[23432] <= r_data[23431];
                
                r_data[23433] <= r_data[23432];
                
                r_data[23434] <= r_data[23433];
                
                r_data[23435] <= r_data[23434];
                
                r_data[23436] <= r_data[23435];
                
                r_data[23437] <= r_data[23436];
                
                r_data[23438] <= r_data[23437];
                
                r_data[23439] <= r_data[23438];
                
                r_data[23440] <= r_data[23439];
                
                r_data[23441] <= r_data[23440];
                
                r_data[23442] <= r_data[23441];
                
                r_data[23443] <= r_data[23442];
                
                r_data[23444] <= r_data[23443];
                
                r_data[23445] <= r_data[23444];
                
                r_data[23446] <= r_data[23445];
                
                r_data[23447] <= r_data[23446];
                
                r_data[23448] <= r_data[23447];
                
                r_data[23449] <= r_data[23448];
                
                r_data[23450] <= r_data[23449];
                
                r_data[23451] <= r_data[23450];
                
                r_data[23452] <= r_data[23451];
                
                r_data[23453] <= r_data[23452];
                
                r_data[23454] <= r_data[23453];
                
                r_data[23455] <= r_data[23454];
                
                r_data[23456] <= r_data[23455];
                
                r_data[23457] <= r_data[23456];
                
                r_data[23458] <= r_data[23457];
                
                r_data[23459] <= r_data[23458];
                
                r_data[23460] <= r_data[23459];
                
                r_data[23461] <= r_data[23460];
                
                r_data[23462] <= r_data[23461];
                
                r_data[23463] <= r_data[23462];
                
                r_data[23464] <= r_data[23463];
                
                r_data[23465] <= r_data[23464];
                
                r_data[23466] <= r_data[23465];
                
                r_data[23467] <= r_data[23466];
                
                r_data[23468] <= r_data[23467];
                
                r_data[23469] <= r_data[23468];
                
                r_data[23470] <= r_data[23469];
                
                r_data[23471] <= r_data[23470];
                
                r_data[23472] <= r_data[23471];
                
                r_data[23473] <= r_data[23472];
                
                r_data[23474] <= r_data[23473];
                
                r_data[23475] <= r_data[23474];
                
                r_data[23476] <= r_data[23475];
                
                r_data[23477] <= r_data[23476];
                
                r_data[23478] <= r_data[23477];
                
                r_data[23479] <= r_data[23478];
                
                r_data[23480] <= r_data[23479];
                
                r_data[23481] <= r_data[23480];
                
                r_data[23482] <= r_data[23481];
                
                r_data[23483] <= r_data[23482];
                
                r_data[23484] <= r_data[23483];
                
                r_data[23485] <= r_data[23484];
                
                r_data[23486] <= r_data[23485];
                
                r_data[23487] <= r_data[23486];
                
                r_data[23488] <= r_data[23487];
                
                r_data[23489] <= r_data[23488];
                
                r_data[23490] <= r_data[23489];
                
                r_data[23491] <= r_data[23490];
                
                r_data[23492] <= r_data[23491];
                
                r_data[23493] <= r_data[23492];
                
                r_data[23494] <= r_data[23493];
                
                r_data[23495] <= r_data[23494];
                
                r_data[23496] <= r_data[23495];
                
                r_data[23497] <= r_data[23496];
                
                r_data[23498] <= r_data[23497];
                
                r_data[23499] <= r_data[23498];
                
                r_data[23500] <= r_data[23499];
                
                r_data[23501] <= r_data[23500];
                
                r_data[23502] <= r_data[23501];
                
                r_data[23503] <= r_data[23502];
                
                r_data[23504] <= r_data[23503];
                
                r_data[23505] <= r_data[23504];
                
                r_data[23506] <= r_data[23505];
                
                r_data[23507] <= r_data[23506];
                
                r_data[23508] <= r_data[23507];
                
                r_data[23509] <= r_data[23508];
                
                r_data[23510] <= r_data[23509];
                
                r_data[23511] <= r_data[23510];
                
                r_data[23512] <= r_data[23511];
                
                r_data[23513] <= r_data[23512];
                
                r_data[23514] <= r_data[23513];
                
                r_data[23515] <= r_data[23514];
                
                r_data[23516] <= r_data[23515];
                
                r_data[23517] <= r_data[23516];
                
                r_data[23518] <= r_data[23517];
                
                r_data[23519] <= r_data[23518];
                
                r_data[23520] <= r_data[23519];
                
                r_data[23521] <= r_data[23520];
                
                r_data[23522] <= r_data[23521];
                
                r_data[23523] <= r_data[23522];
                
                r_data[23524] <= r_data[23523];
                
                r_data[23525] <= r_data[23524];
                
                r_data[23526] <= r_data[23525];
                
                r_data[23527] <= r_data[23526];
                
                r_data[23528] <= r_data[23527];
                
                r_data[23529] <= r_data[23528];
                
                r_data[23530] <= r_data[23529];
                
                r_data[23531] <= r_data[23530];
                
                r_data[23532] <= r_data[23531];
                
                r_data[23533] <= r_data[23532];
                
                r_data[23534] <= r_data[23533];
                
                r_data[23535] <= r_data[23534];
                
                r_data[23536] <= r_data[23535];
                
                r_data[23537] <= r_data[23536];
                
                r_data[23538] <= r_data[23537];
                
                r_data[23539] <= r_data[23538];
                
                r_data[23540] <= r_data[23539];
                
                r_data[23541] <= r_data[23540];
                
                r_data[23542] <= r_data[23541];
                
                r_data[23543] <= r_data[23542];
                
                r_data[23544] <= r_data[23543];
                
                r_data[23545] <= r_data[23544];
                
                r_data[23546] <= r_data[23545];
                
                r_data[23547] <= r_data[23546];
                
                r_data[23548] <= r_data[23547];
                
                r_data[23549] <= r_data[23548];
                
                r_data[23550] <= r_data[23549];
                
                r_data[23551] <= r_data[23550];
                
                r_data[23552] <= r_data[23551];
                
                r_data[23553] <= r_data[23552];
                
                r_data[23554] <= r_data[23553];
                
                r_data[23555] <= r_data[23554];
                
                r_data[23556] <= r_data[23555];
                
                r_data[23557] <= r_data[23556];
                
                r_data[23558] <= r_data[23557];
                
                r_data[23559] <= r_data[23558];
                
                r_data[23560] <= r_data[23559];
                
                r_data[23561] <= r_data[23560];
                
                r_data[23562] <= r_data[23561];
                
                r_data[23563] <= r_data[23562];
                
                r_data[23564] <= r_data[23563];
                
                r_data[23565] <= r_data[23564];
                
                r_data[23566] <= r_data[23565];
                
                r_data[23567] <= r_data[23566];
                
                r_data[23568] <= r_data[23567];
                
                r_data[23569] <= r_data[23568];
                
                r_data[23570] <= r_data[23569];
                
                r_data[23571] <= r_data[23570];
                
                r_data[23572] <= r_data[23571];
                
                r_data[23573] <= r_data[23572];
                
                r_data[23574] <= r_data[23573];
                
                r_data[23575] <= r_data[23574];
                
                r_data[23576] <= r_data[23575];
                
                r_data[23577] <= r_data[23576];
                
                r_data[23578] <= r_data[23577];
                
                r_data[23579] <= r_data[23578];
                
                r_data[23580] <= r_data[23579];
                
                r_data[23581] <= r_data[23580];
                
                r_data[23582] <= r_data[23581];
                
                r_data[23583] <= r_data[23582];
                
                r_data[23584] <= r_data[23583];
                
                r_data[23585] <= r_data[23584];
                
                r_data[23586] <= r_data[23585];
                
                r_data[23587] <= r_data[23586];
                
                r_data[23588] <= r_data[23587];
                
                r_data[23589] <= r_data[23588];
                
                r_data[23590] <= r_data[23589];
                
                r_data[23591] <= r_data[23590];
                
                r_data[23592] <= r_data[23591];
                
                r_data[23593] <= r_data[23592];
                
                r_data[23594] <= r_data[23593];
                
                r_data[23595] <= r_data[23594];
                
                r_data[23596] <= r_data[23595];
                
                r_data[23597] <= r_data[23596];
                
                r_data[23598] <= r_data[23597];
                
                r_data[23599] <= r_data[23598];
                
                r_data[23600] <= r_data[23599];
                
                r_data[23601] <= r_data[23600];
                
                r_data[23602] <= r_data[23601];
                
                r_data[23603] <= r_data[23602];
                
                r_data[23604] <= r_data[23603];
                
                r_data[23605] <= r_data[23604];
                
                r_data[23606] <= r_data[23605];
                
                r_data[23607] <= r_data[23606];
                
                r_data[23608] <= r_data[23607];
                
                r_data[23609] <= r_data[23608];
                
                r_data[23610] <= r_data[23609];
                
                r_data[23611] <= r_data[23610];
                
                r_data[23612] <= r_data[23611];
                
                r_data[23613] <= r_data[23612];
                
                r_data[23614] <= r_data[23613];
                
                r_data[23615] <= r_data[23614];
                
                r_data[23616] <= r_data[23615];
                
                r_data[23617] <= r_data[23616];
                
                r_data[23618] <= r_data[23617];
                
                r_data[23619] <= r_data[23618];
                
                r_data[23620] <= r_data[23619];
                
                r_data[23621] <= r_data[23620];
                
                r_data[23622] <= r_data[23621];
                
                r_data[23623] <= r_data[23622];
                
                r_data[23624] <= r_data[23623];
                
                r_data[23625] <= r_data[23624];
                
                r_data[23626] <= r_data[23625];
                
                r_data[23627] <= r_data[23626];
                
                r_data[23628] <= r_data[23627];
                
                r_data[23629] <= r_data[23628];
                
                r_data[23630] <= r_data[23629];
                
                r_data[23631] <= r_data[23630];
                
                r_data[23632] <= r_data[23631];
                
                r_data[23633] <= r_data[23632];
                
                r_data[23634] <= r_data[23633];
                
                r_data[23635] <= r_data[23634];
                
                r_data[23636] <= r_data[23635];
                
                r_data[23637] <= r_data[23636];
                
                r_data[23638] <= r_data[23637];
                
                r_data[23639] <= r_data[23638];
                
                r_data[23640] <= r_data[23639];
                
                r_data[23641] <= r_data[23640];
                
                r_data[23642] <= r_data[23641];
                
                r_data[23643] <= r_data[23642];
                
                r_data[23644] <= r_data[23643];
                
                r_data[23645] <= r_data[23644];
                
                r_data[23646] <= r_data[23645];
                
                r_data[23647] <= r_data[23646];
                
                r_data[23648] <= r_data[23647];
                
                r_data[23649] <= r_data[23648];
                
                r_data[23650] <= r_data[23649];
                
                r_data[23651] <= r_data[23650];
                
                r_data[23652] <= r_data[23651];
                
                r_data[23653] <= r_data[23652];
                
                r_data[23654] <= r_data[23653];
                
                r_data[23655] <= r_data[23654];
                
                r_data[23656] <= r_data[23655];
                
                r_data[23657] <= r_data[23656];
                
                r_data[23658] <= r_data[23657];
                
                r_data[23659] <= r_data[23658];
                
                r_data[23660] <= r_data[23659];
                
                r_data[23661] <= r_data[23660];
                
                r_data[23662] <= r_data[23661];
                
                r_data[23663] <= r_data[23662];
                
                r_data[23664] <= r_data[23663];
                
                r_data[23665] <= r_data[23664];
                
                r_data[23666] <= r_data[23665];
                
                r_data[23667] <= r_data[23666];
                
                r_data[23668] <= r_data[23667];
                
                r_data[23669] <= r_data[23668];
                
                r_data[23670] <= r_data[23669];
                
                r_data[23671] <= r_data[23670];
                
                r_data[23672] <= r_data[23671];
                
                r_data[23673] <= r_data[23672];
                
                r_data[23674] <= r_data[23673];
                
                r_data[23675] <= r_data[23674];
                
                r_data[23676] <= r_data[23675];
                
                r_data[23677] <= r_data[23676];
                
                r_data[23678] <= r_data[23677];
                
                r_data[23679] <= r_data[23678];
                
                r_data[23680] <= r_data[23679];
                
                r_data[23681] <= r_data[23680];
                
                r_data[23682] <= r_data[23681];
                
                r_data[23683] <= r_data[23682];
                
                r_data[23684] <= r_data[23683];
                
                r_data[23685] <= r_data[23684];
                
                r_data[23686] <= r_data[23685];
                
                r_data[23687] <= r_data[23686];
                
                r_data[23688] <= r_data[23687];
                
                r_data[23689] <= r_data[23688];
                
                r_data[23690] <= r_data[23689];
                
                r_data[23691] <= r_data[23690];
                
                r_data[23692] <= r_data[23691];
                
                r_data[23693] <= r_data[23692];
                
                r_data[23694] <= r_data[23693];
                
                r_data[23695] <= r_data[23694];
                
                r_data[23696] <= r_data[23695];
                
                r_data[23697] <= r_data[23696];
                
                r_data[23698] <= r_data[23697];
                
                r_data[23699] <= r_data[23698];
                
                r_data[23700] <= r_data[23699];
                
                r_data[23701] <= r_data[23700];
                
                r_data[23702] <= r_data[23701];
                
                r_data[23703] <= r_data[23702];
                
                r_data[23704] <= r_data[23703];
                
                r_data[23705] <= r_data[23704];
                
                r_data[23706] <= r_data[23705];
                
                r_data[23707] <= r_data[23706];
                
                r_data[23708] <= r_data[23707];
                
                r_data[23709] <= r_data[23708];
                
                r_data[23710] <= r_data[23709];
                
                r_data[23711] <= r_data[23710];
                
                r_data[23712] <= r_data[23711];
                
                r_data[23713] <= r_data[23712];
                
                r_data[23714] <= r_data[23713];
                
                r_data[23715] <= r_data[23714];
                
                r_data[23716] <= r_data[23715];
                
                r_data[23717] <= r_data[23716];
                
                r_data[23718] <= r_data[23717];
                
                r_data[23719] <= r_data[23718];
                
                r_data[23720] <= r_data[23719];
                
                r_data[23721] <= r_data[23720];
                
                r_data[23722] <= r_data[23721];
                
                r_data[23723] <= r_data[23722];
                
                r_data[23724] <= r_data[23723];
                
                r_data[23725] <= r_data[23724];
                
                r_data[23726] <= r_data[23725];
                
                r_data[23727] <= r_data[23726];
                
                r_data[23728] <= r_data[23727];
                
                r_data[23729] <= r_data[23728];
                
                r_data[23730] <= r_data[23729];
                
                r_data[23731] <= r_data[23730];
                
                r_data[23732] <= r_data[23731];
                
                r_data[23733] <= r_data[23732];
                
                r_data[23734] <= r_data[23733];
                
                r_data[23735] <= r_data[23734];
                
                r_data[23736] <= r_data[23735];
                
                r_data[23737] <= r_data[23736];
                
                r_data[23738] <= r_data[23737];
                
                r_data[23739] <= r_data[23738];
                
                r_data[23740] <= r_data[23739];
                
                r_data[23741] <= r_data[23740];
                
                r_data[23742] <= r_data[23741];
                
                r_data[23743] <= r_data[23742];
                
                r_data[23744] <= r_data[23743];
                
                r_data[23745] <= r_data[23744];
                
                r_data[23746] <= r_data[23745];
                
                r_data[23747] <= r_data[23746];
                
                r_data[23748] <= r_data[23747];
                
                r_data[23749] <= r_data[23748];
                
                r_data[23750] <= r_data[23749];
                
                r_data[23751] <= r_data[23750];
                
                r_data[23752] <= r_data[23751];
                
                r_data[23753] <= r_data[23752];
                
                r_data[23754] <= r_data[23753];
                
                r_data[23755] <= r_data[23754];
                
                r_data[23756] <= r_data[23755];
                
                r_data[23757] <= r_data[23756];
                
                r_data[23758] <= r_data[23757];
                
                r_data[23759] <= r_data[23758];
                
                r_data[23760] <= r_data[23759];
                
                r_data[23761] <= r_data[23760];
                
                r_data[23762] <= r_data[23761];
                
                r_data[23763] <= r_data[23762];
                
                r_data[23764] <= r_data[23763];
                
                r_data[23765] <= r_data[23764];
                
                r_data[23766] <= r_data[23765];
                
                r_data[23767] <= r_data[23766];
                
                r_data[23768] <= r_data[23767];
                
                r_data[23769] <= r_data[23768];
                
                r_data[23770] <= r_data[23769];
                
                r_data[23771] <= r_data[23770];
                
                r_data[23772] <= r_data[23771];
                
                r_data[23773] <= r_data[23772];
                
                r_data[23774] <= r_data[23773];
                
                r_data[23775] <= r_data[23774];
                
                r_data[23776] <= r_data[23775];
                
                r_data[23777] <= r_data[23776];
                
                r_data[23778] <= r_data[23777];
                
                r_data[23779] <= r_data[23778];
                
                r_data[23780] <= r_data[23779];
                
                r_data[23781] <= r_data[23780];
                
                r_data[23782] <= r_data[23781];
                
                r_data[23783] <= r_data[23782];
                
                r_data[23784] <= r_data[23783];
                
                r_data[23785] <= r_data[23784];
                
                r_data[23786] <= r_data[23785];
                
                r_data[23787] <= r_data[23786];
                
                r_data[23788] <= r_data[23787];
                
                r_data[23789] <= r_data[23788];
                
                r_data[23790] <= r_data[23789];
                
                r_data[23791] <= r_data[23790];
                
                r_data[23792] <= r_data[23791];
                
                r_data[23793] <= r_data[23792];
                
                r_data[23794] <= r_data[23793];
                
                r_data[23795] <= r_data[23794];
                
                r_data[23796] <= r_data[23795];
                
                r_data[23797] <= r_data[23796];
                
                r_data[23798] <= r_data[23797];
                
                r_data[23799] <= r_data[23798];
                
                r_data[23800] <= r_data[23799];
                
                r_data[23801] <= r_data[23800];
                
                r_data[23802] <= r_data[23801];
                
                r_data[23803] <= r_data[23802];
                
                r_data[23804] <= r_data[23803];
                
                r_data[23805] <= r_data[23804];
                
                r_data[23806] <= r_data[23805];
                
                r_data[23807] <= r_data[23806];
                
                r_data[23808] <= r_data[23807];
                
                r_data[23809] <= r_data[23808];
                
                r_data[23810] <= r_data[23809];
                
                r_data[23811] <= r_data[23810];
                
                r_data[23812] <= r_data[23811];
                
                r_data[23813] <= r_data[23812];
                
                r_data[23814] <= r_data[23813];
                
                r_data[23815] <= r_data[23814];
                
                r_data[23816] <= r_data[23815];
                
                r_data[23817] <= r_data[23816];
                
                r_data[23818] <= r_data[23817];
                
                r_data[23819] <= r_data[23818];
                
                r_data[23820] <= r_data[23819];
                
                r_data[23821] <= r_data[23820];
                
                r_data[23822] <= r_data[23821];
                
                r_data[23823] <= r_data[23822];
                
                r_data[23824] <= r_data[23823];
                
                r_data[23825] <= r_data[23824];
                
                r_data[23826] <= r_data[23825];
                
                r_data[23827] <= r_data[23826];
                
                r_data[23828] <= r_data[23827];
                
                r_data[23829] <= r_data[23828];
                
                r_data[23830] <= r_data[23829];
                
                r_data[23831] <= r_data[23830];
                
                r_data[23832] <= r_data[23831];
                
                r_data[23833] <= r_data[23832];
                
                r_data[23834] <= r_data[23833];
                
                r_data[23835] <= r_data[23834];
                
                r_data[23836] <= r_data[23835];
                
                r_data[23837] <= r_data[23836];
                
                r_data[23838] <= r_data[23837];
                
                r_data[23839] <= r_data[23838];
                
                r_data[23840] <= r_data[23839];
                
                r_data[23841] <= r_data[23840];
                
                r_data[23842] <= r_data[23841];
                
                r_data[23843] <= r_data[23842];
                
                r_data[23844] <= r_data[23843];
                
                r_data[23845] <= r_data[23844];
                
                r_data[23846] <= r_data[23845];
                
                r_data[23847] <= r_data[23846];
                
                r_data[23848] <= r_data[23847];
                
                r_data[23849] <= r_data[23848];
                
                r_data[23850] <= r_data[23849];
                
                r_data[23851] <= r_data[23850];
                
                r_data[23852] <= r_data[23851];
                
                r_data[23853] <= r_data[23852];
                
                r_data[23854] <= r_data[23853];
                
                r_data[23855] <= r_data[23854];
                
                r_data[23856] <= r_data[23855];
                
                r_data[23857] <= r_data[23856];
                
                r_data[23858] <= r_data[23857];
                
                r_data[23859] <= r_data[23858];
                
                r_data[23860] <= r_data[23859];
                
                r_data[23861] <= r_data[23860];
                
                r_data[23862] <= r_data[23861];
                
                r_data[23863] <= r_data[23862];
                
                r_data[23864] <= r_data[23863];
                
                r_data[23865] <= r_data[23864];
                
                r_data[23866] <= r_data[23865];
                
                r_data[23867] <= r_data[23866];
                
                r_data[23868] <= r_data[23867];
                
                r_data[23869] <= r_data[23868];
                
                r_data[23870] <= r_data[23869];
                
                r_data[23871] <= r_data[23870];
                
                r_data[23872] <= r_data[23871];
                
                r_data[23873] <= r_data[23872];
                
                r_data[23874] <= r_data[23873];
                
                r_data[23875] <= r_data[23874];
                
                r_data[23876] <= r_data[23875];
                
                r_data[23877] <= r_data[23876];
                
                r_data[23878] <= r_data[23877];
                
                r_data[23879] <= r_data[23878];
                
                r_data[23880] <= r_data[23879];
                
                r_data[23881] <= r_data[23880];
                
                r_data[23882] <= r_data[23881];
                
                r_data[23883] <= r_data[23882];
                
                r_data[23884] <= r_data[23883];
                
                r_data[23885] <= r_data[23884];
                
                r_data[23886] <= r_data[23885];
                
                r_data[23887] <= r_data[23886];
                
                r_data[23888] <= r_data[23887];
                
                r_data[23889] <= r_data[23888];
                
                r_data[23890] <= r_data[23889];
                
                r_data[23891] <= r_data[23890];
                
                r_data[23892] <= r_data[23891];
                
                r_data[23893] <= r_data[23892];
                
                r_data[23894] <= r_data[23893];
                
                r_data[23895] <= r_data[23894];
                
                r_data[23896] <= r_data[23895];
                
                r_data[23897] <= r_data[23896];
                
                r_data[23898] <= r_data[23897];
                
                r_data[23899] <= r_data[23898];
                
                r_data[23900] <= r_data[23899];
                
                r_data[23901] <= r_data[23900];
                
                r_data[23902] <= r_data[23901];
                
                r_data[23903] <= r_data[23902];
                
                r_data[23904] <= r_data[23903];
                
                r_data[23905] <= r_data[23904];
                
                r_data[23906] <= r_data[23905];
                
                r_data[23907] <= r_data[23906];
                
                r_data[23908] <= r_data[23907];
                
                r_data[23909] <= r_data[23908];
                
                r_data[23910] <= r_data[23909];
                
                r_data[23911] <= r_data[23910];
                
                r_data[23912] <= r_data[23911];
                
                r_data[23913] <= r_data[23912];
                
                r_data[23914] <= r_data[23913];
                
                r_data[23915] <= r_data[23914];
                
                r_data[23916] <= r_data[23915];
                
                r_data[23917] <= r_data[23916];
                
                r_data[23918] <= r_data[23917];
                
                r_data[23919] <= r_data[23918];
                
                r_data[23920] <= r_data[23919];
                
                r_data[23921] <= r_data[23920];
                
                r_data[23922] <= r_data[23921];
                
                r_data[23923] <= r_data[23922];
                
                r_data[23924] <= r_data[23923];
                
                r_data[23925] <= r_data[23924];
                
                r_data[23926] <= r_data[23925];
                
                r_data[23927] <= r_data[23926];
                
                r_data[23928] <= r_data[23927];
                
                r_data[23929] <= r_data[23928];
                
                r_data[23930] <= r_data[23929];
                
                r_data[23931] <= r_data[23930];
                
                r_data[23932] <= r_data[23931];
                
                r_data[23933] <= r_data[23932];
                
                r_data[23934] <= r_data[23933];
                
                r_data[23935] <= r_data[23934];
                
                r_data[23936] <= r_data[23935];
                
                r_data[23937] <= r_data[23936];
                
                r_data[23938] <= r_data[23937];
                
                r_data[23939] <= r_data[23938];
                
                r_data[23940] <= r_data[23939];
                
                r_data[23941] <= r_data[23940];
                
                r_data[23942] <= r_data[23941];
                
                r_data[23943] <= r_data[23942];
                
                r_data[23944] <= r_data[23943];
                
                r_data[23945] <= r_data[23944];
                
                r_data[23946] <= r_data[23945];
                
                r_data[23947] <= r_data[23946];
                
                r_data[23948] <= r_data[23947];
                
                r_data[23949] <= r_data[23948];
                
                r_data[23950] <= r_data[23949];
                
                r_data[23951] <= r_data[23950];
                
                r_data[23952] <= r_data[23951];
                
                r_data[23953] <= r_data[23952];
                
                r_data[23954] <= r_data[23953];
                
                r_data[23955] <= r_data[23954];
                
                r_data[23956] <= r_data[23955];
                
                r_data[23957] <= r_data[23956];
                
                r_data[23958] <= r_data[23957];
                
                r_data[23959] <= r_data[23958];
                
                r_data[23960] <= r_data[23959];
                
                r_data[23961] <= r_data[23960];
                
                r_data[23962] <= r_data[23961];
                
                r_data[23963] <= r_data[23962];
                
                r_data[23964] <= r_data[23963];
                
                r_data[23965] <= r_data[23964];
                
                r_data[23966] <= r_data[23965];
                
                r_data[23967] <= r_data[23966];
                
                r_data[23968] <= r_data[23967];
                
                r_data[23969] <= r_data[23968];
                
                r_data[23970] <= r_data[23969];
                
                r_data[23971] <= r_data[23970];
                
                r_data[23972] <= r_data[23971];
                
                r_data[23973] <= r_data[23972];
                
                r_data[23974] <= r_data[23973];
                
                r_data[23975] <= r_data[23974];
                
                r_data[23976] <= r_data[23975];
                
                r_data[23977] <= r_data[23976];
                
                r_data[23978] <= r_data[23977];
                
                r_data[23979] <= r_data[23978];
                
                r_data[23980] <= r_data[23979];
                
                r_data[23981] <= r_data[23980];
                
                r_data[23982] <= r_data[23981];
                
                r_data[23983] <= r_data[23982];
                
                r_data[23984] <= r_data[23983];
                
                r_data[23985] <= r_data[23984];
                
                r_data[23986] <= r_data[23985];
                
                r_data[23987] <= r_data[23986];
                
                r_data[23988] <= r_data[23987];
                
                r_data[23989] <= r_data[23988];
                
                r_data[23990] <= r_data[23989];
                
                r_data[23991] <= r_data[23990];
                
                r_data[23992] <= r_data[23991];
                
                r_data[23993] <= r_data[23992];
                
                r_data[23994] <= r_data[23993];
                
                r_data[23995] <= r_data[23994];
                
                r_data[23996] <= r_data[23995];
                
                r_data[23997] <= r_data[23996];
                
                r_data[23998] <= r_data[23997];
                
                r_data[23999] <= r_data[23998];
                
                r_data[24000] <= r_data[23999];
                
                r_data[24001] <= r_data[24000];
                
                r_data[24002] <= r_data[24001];
                
                r_data[24003] <= r_data[24002];
                
                r_data[24004] <= r_data[24003];
                
                r_data[24005] <= r_data[24004];
                
                r_data[24006] <= r_data[24005];
                
                r_data[24007] <= r_data[24006];
                
                r_data[24008] <= r_data[24007];
                
                r_data[24009] <= r_data[24008];
                
                r_data[24010] <= r_data[24009];
                
                r_data[24011] <= r_data[24010];
                
                r_data[24012] <= r_data[24011];
                
                r_data[24013] <= r_data[24012];
                
                r_data[24014] <= r_data[24013];
                
                r_data[24015] <= r_data[24014];
                
                r_data[24016] <= r_data[24015];
                
                r_data[24017] <= r_data[24016];
                
                r_data[24018] <= r_data[24017];
                
                r_data[24019] <= r_data[24018];
                
                r_data[24020] <= r_data[24019];
                
                r_data[24021] <= r_data[24020];
                
                r_data[24022] <= r_data[24021];
                
                r_data[24023] <= r_data[24022];
                
                r_data[24024] <= r_data[24023];
                
                r_data[24025] <= r_data[24024];
                
                r_data[24026] <= r_data[24025];
                
                r_data[24027] <= r_data[24026];
                
                r_data[24028] <= r_data[24027];
                
                r_data[24029] <= r_data[24028];
                
                r_data[24030] <= r_data[24029];
                
                r_data[24031] <= r_data[24030];
                
                r_data[24032] <= r_data[24031];
                
                r_data[24033] <= r_data[24032];
                
                r_data[24034] <= r_data[24033];
                
                r_data[24035] <= r_data[24034];
                
                r_data[24036] <= r_data[24035];
                
                r_data[24037] <= r_data[24036];
                
                r_data[24038] <= r_data[24037];
                
                r_data[24039] <= r_data[24038];
                
                r_data[24040] <= r_data[24039];
                
                r_data[24041] <= r_data[24040];
                
                r_data[24042] <= r_data[24041];
                
                r_data[24043] <= r_data[24042];
                
                r_data[24044] <= r_data[24043];
                
                r_data[24045] <= r_data[24044];
                
                r_data[24046] <= r_data[24045];
                
                r_data[24047] <= r_data[24046];
                
                r_data[24048] <= r_data[24047];
                
                r_data[24049] <= r_data[24048];
                
                r_data[24050] <= r_data[24049];
                
                r_data[24051] <= r_data[24050];
                
                r_data[24052] <= r_data[24051];
                
                r_data[24053] <= r_data[24052];
                
                r_data[24054] <= r_data[24053];
                
                r_data[24055] <= r_data[24054];
                
                r_data[24056] <= r_data[24055];
                
                r_data[24057] <= r_data[24056];
                
                r_data[24058] <= r_data[24057];
                
                r_data[24059] <= r_data[24058];
                
                r_data[24060] <= r_data[24059];
                
                r_data[24061] <= r_data[24060];
                
                r_data[24062] <= r_data[24061];
                
                r_data[24063] <= r_data[24062];
                
                r_data[24064] <= r_data[24063];
                
                r_data[24065] <= r_data[24064];
                
                r_data[24066] <= r_data[24065];
                
                r_data[24067] <= r_data[24066];
                
                r_data[24068] <= r_data[24067];
                
                r_data[24069] <= r_data[24068];
                
                r_data[24070] <= r_data[24069];
                
                r_data[24071] <= r_data[24070];
                
                r_data[24072] <= r_data[24071];
                
                r_data[24073] <= r_data[24072];
                
                r_data[24074] <= r_data[24073];
                
                r_data[24075] <= r_data[24074];
                
                r_data[24076] <= r_data[24075];
                
                r_data[24077] <= r_data[24076];
                
                r_data[24078] <= r_data[24077];
                
                r_data[24079] <= r_data[24078];
                
                r_data[24080] <= r_data[24079];
                
                r_data[24081] <= r_data[24080];
                
                r_data[24082] <= r_data[24081];
                
                r_data[24083] <= r_data[24082];
                
                r_data[24084] <= r_data[24083];
                
                r_data[24085] <= r_data[24084];
                
                r_data[24086] <= r_data[24085];
                
                r_data[24087] <= r_data[24086];
                
                r_data[24088] <= r_data[24087];
                
                r_data[24089] <= r_data[24088];
                
                r_data[24090] <= r_data[24089];
                
                r_data[24091] <= r_data[24090];
                
                r_data[24092] <= r_data[24091];
                
                r_data[24093] <= r_data[24092];
                
                r_data[24094] <= r_data[24093];
                
                r_data[24095] <= r_data[24094];
                
                r_data[24096] <= r_data[24095];
                
                r_data[24097] <= r_data[24096];
                
                r_data[24098] <= r_data[24097];
                
                r_data[24099] <= r_data[24098];
                
                r_data[24100] <= r_data[24099];
                
                r_data[24101] <= r_data[24100];
                
                r_data[24102] <= r_data[24101];
                
                r_data[24103] <= r_data[24102];
                
                r_data[24104] <= r_data[24103];
                
                r_data[24105] <= r_data[24104];
                
                r_data[24106] <= r_data[24105];
                
                r_data[24107] <= r_data[24106];
                
                r_data[24108] <= r_data[24107];
                
                r_data[24109] <= r_data[24108];
                
                r_data[24110] <= r_data[24109];
                
                r_data[24111] <= r_data[24110];
                
                r_data[24112] <= r_data[24111];
                
                r_data[24113] <= r_data[24112];
                
                r_data[24114] <= r_data[24113];
                
                r_data[24115] <= r_data[24114];
                
                r_data[24116] <= r_data[24115];
                
                r_data[24117] <= r_data[24116];
                
                r_data[24118] <= r_data[24117];
                
                r_data[24119] <= r_data[24118];
                
                r_data[24120] <= r_data[24119];
                
                r_data[24121] <= r_data[24120];
                
                r_data[24122] <= r_data[24121];
                
                r_data[24123] <= r_data[24122];
                
                r_data[24124] <= r_data[24123];
                
                r_data[24125] <= r_data[24124];
                
                r_data[24126] <= r_data[24125];
                
                r_data[24127] <= r_data[24126];
                
                r_data[24128] <= r_data[24127];
                
                r_data[24129] <= r_data[24128];
                
                r_data[24130] <= r_data[24129];
                
                r_data[24131] <= r_data[24130];
                
                r_data[24132] <= r_data[24131];
                
                r_data[24133] <= r_data[24132];
                
                r_data[24134] <= r_data[24133];
                
                r_data[24135] <= r_data[24134];
                
                r_data[24136] <= r_data[24135];
                
                r_data[24137] <= r_data[24136];
                
                r_data[24138] <= r_data[24137];
                
                r_data[24139] <= r_data[24138];
                
                r_data[24140] <= r_data[24139];
                
                r_data[24141] <= r_data[24140];
                
                r_data[24142] <= r_data[24141];
                
                r_data[24143] <= r_data[24142];
                
                r_data[24144] <= r_data[24143];
                
                r_data[24145] <= r_data[24144];
                
                r_data[24146] <= r_data[24145];
                
                r_data[24147] <= r_data[24146];
                
                r_data[24148] <= r_data[24147];
                
                r_data[24149] <= r_data[24148];
                
                r_data[24150] <= r_data[24149];
                
                r_data[24151] <= r_data[24150];
                
                r_data[24152] <= r_data[24151];
                
                r_data[24153] <= r_data[24152];
                
                r_data[24154] <= r_data[24153];
                
                r_data[24155] <= r_data[24154];
                
                r_data[24156] <= r_data[24155];
                
                r_data[24157] <= r_data[24156];
                
                r_data[24158] <= r_data[24157];
                
                r_data[24159] <= r_data[24158];
                
                r_data[24160] <= r_data[24159];
                
                r_data[24161] <= r_data[24160];
                
                r_data[24162] <= r_data[24161];
                
                r_data[24163] <= r_data[24162];
                
                r_data[24164] <= r_data[24163];
                
                r_data[24165] <= r_data[24164];
                
                r_data[24166] <= r_data[24165];
                
                r_data[24167] <= r_data[24166];
                
                r_data[24168] <= r_data[24167];
                
                r_data[24169] <= r_data[24168];
                
                r_data[24170] <= r_data[24169];
                
                r_data[24171] <= r_data[24170];
                
                r_data[24172] <= r_data[24171];
                
                r_data[24173] <= r_data[24172];
                
                r_data[24174] <= r_data[24173];
                
                r_data[24175] <= r_data[24174];
                
                r_data[24176] <= r_data[24175];
                
                r_data[24177] <= r_data[24176];
                
                r_data[24178] <= r_data[24177];
                
                r_data[24179] <= r_data[24178];
                
                r_data[24180] <= r_data[24179];
                
                r_data[24181] <= r_data[24180];
                
                r_data[24182] <= r_data[24181];
                
                r_data[24183] <= r_data[24182];
                
                r_data[24184] <= r_data[24183];
                
                r_data[24185] <= r_data[24184];
                
                r_data[24186] <= r_data[24185];
                
                r_data[24187] <= r_data[24186];
                
                r_data[24188] <= r_data[24187];
                
                r_data[24189] <= r_data[24188];
                
                r_data[24190] <= r_data[24189];
                
                r_data[24191] <= r_data[24190];
                
                r_data[24192] <= r_data[24191];
                
                r_data[24193] <= r_data[24192];
                
                r_data[24194] <= r_data[24193];
                
                r_data[24195] <= r_data[24194];
                
                r_data[24196] <= r_data[24195];
                
                r_data[24197] <= r_data[24196];
                
                r_data[24198] <= r_data[24197];
                
                r_data[24199] <= r_data[24198];
                
                r_data[24200] <= r_data[24199];
                
                r_data[24201] <= r_data[24200];
                
                r_data[24202] <= r_data[24201];
                
                r_data[24203] <= r_data[24202];
                
                r_data[24204] <= r_data[24203];
                
                r_data[24205] <= r_data[24204];
                
                r_data[24206] <= r_data[24205];
                
                r_data[24207] <= r_data[24206];
                
                r_data[24208] <= r_data[24207];
                
                r_data[24209] <= r_data[24208];
                
                r_data[24210] <= r_data[24209];
                
                r_data[24211] <= r_data[24210];
                
                r_data[24212] <= r_data[24211];
                
                r_data[24213] <= r_data[24212];
                
                r_data[24214] <= r_data[24213];
                
                r_data[24215] <= r_data[24214];
                
                r_data[24216] <= r_data[24215];
                
                r_data[24217] <= r_data[24216];
                
                r_data[24218] <= r_data[24217];
                
                r_data[24219] <= r_data[24218];
                
                r_data[24220] <= r_data[24219];
                
                r_data[24221] <= r_data[24220];
                
                r_data[24222] <= r_data[24221];
                
                r_data[24223] <= r_data[24222];
                
                r_data[24224] <= r_data[24223];
                
                r_data[24225] <= r_data[24224];
                
                r_data[24226] <= r_data[24225];
                
                r_data[24227] <= r_data[24226];
                
                r_data[24228] <= r_data[24227];
                
                r_data[24229] <= r_data[24228];
                
                r_data[24230] <= r_data[24229];
                
                r_data[24231] <= r_data[24230];
                
                r_data[24232] <= r_data[24231];
                
                r_data[24233] <= r_data[24232];
                
                r_data[24234] <= r_data[24233];
                
                r_data[24235] <= r_data[24234];
                
                r_data[24236] <= r_data[24235];
                
                r_data[24237] <= r_data[24236];
                
                r_data[24238] <= r_data[24237];
                
                r_data[24239] <= r_data[24238];
                
                r_data[24240] <= r_data[24239];
                
                r_data[24241] <= r_data[24240];
                
                r_data[24242] <= r_data[24241];
                
                r_data[24243] <= r_data[24242];
                
                r_data[24244] <= r_data[24243];
                
                r_data[24245] <= r_data[24244];
                
                r_data[24246] <= r_data[24245];
                
                r_data[24247] <= r_data[24246];
                
                r_data[24248] <= r_data[24247];
                
                r_data[24249] <= r_data[24248];
                
                r_data[24250] <= r_data[24249];
                
                r_data[24251] <= r_data[24250];
                
                r_data[24252] <= r_data[24251];
                
                r_data[24253] <= r_data[24252];
                
                r_data[24254] <= r_data[24253];
                
                r_data[24255] <= r_data[24254];
                
                r_data[24256] <= r_data[24255];
                
                r_data[24257] <= r_data[24256];
                
                r_data[24258] <= r_data[24257];
                
                r_data[24259] <= r_data[24258];
                
                r_data[24260] <= r_data[24259];
                
                r_data[24261] <= r_data[24260];
                
                r_data[24262] <= r_data[24261];
                
                r_data[24263] <= r_data[24262];
                
                r_data[24264] <= r_data[24263];
                
                r_data[24265] <= r_data[24264];
                
                r_data[24266] <= r_data[24265];
                
                r_data[24267] <= r_data[24266];
                
                r_data[24268] <= r_data[24267];
                
                r_data[24269] <= r_data[24268];
                
                r_data[24270] <= r_data[24269];
                
                r_data[24271] <= r_data[24270];
                
                r_data[24272] <= r_data[24271];
                
                r_data[24273] <= r_data[24272];
                
                r_data[24274] <= r_data[24273];
                
                r_data[24275] <= r_data[24274];
                
                r_data[24276] <= r_data[24275];
                
                r_data[24277] <= r_data[24276];
                
                r_data[24278] <= r_data[24277];
                
                r_data[24279] <= r_data[24278];
                
                r_data[24280] <= r_data[24279];
                
                r_data[24281] <= r_data[24280];
                
                r_data[24282] <= r_data[24281];
                
                r_data[24283] <= r_data[24282];
                
                r_data[24284] <= r_data[24283];
                
                r_data[24285] <= r_data[24284];
                
                r_data[24286] <= r_data[24285];
                
                r_data[24287] <= r_data[24286];
                
                r_data[24288] <= r_data[24287];
                
                r_data[24289] <= r_data[24288];
                
                r_data[24290] <= r_data[24289];
                
                r_data[24291] <= r_data[24290];
                
                r_data[24292] <= r_data[24291];
                
                r_data[24293] <= r_data[24292];
                
                r_data[24294] <= r_data[24293];
                
                r_data[24295] <= r_data[24294];
                
                r_data[24296] <= r_data[24295];
                
                r_data[24297] <= r_data[24296];
                
                r_data[24298] <= r_data[24297];
                
                r_data[24299] <= r_data[24298];
                
                r_data[24300] <= r_data[24299];
                
                r_data[24301] <= r_data[24300];
                
                r_data[24302] <= r_data[24301];
                
                r_data[24303] <= r_data[24302];
                
                r_data[24304] <= r_data[24303];
                
                r_data[24305] <= r_data[24304];
                
                r_data[24306] <= r_data[24305];
                
                r_data[24307] <= r_data[24306];
                
                r_data[24308] <= r_data[24307];
                
                r_data[24309] <= r_data[24308];
                
                r_data[24310] <= r_data[24309];
                
                r_data[24311] <= r_data[24310];
                
                r_data[24312] <= r_data[24311];
                
                r_data[24313] <= r_data[24312];
                
                r_data[24314] <= r_data[24313];
                
                r_data[24315] <= r_data[24314];
                
                r_data[24316] <= r_data[24315];
                
                r_data[24317] <= r_data[24316];
                
                r_data[24318] <= r_data[24317];
                
                r_data[24319] <= r_data[24318];
                
                r_data[24320] <= r_data[24319];
                
                r_data[24321] <= r_data[24320];
                
                r_data[24322] <= r_data[24321];
                
                r_data[24323] <= r_data[24322];
                
                r_data[24324] <= r_data[24323];
                
                r_data[24325] <= r_data[24324];
                
                r_data[24326] <= r_data[24325];
                
                r_data[24327] <= r_data[24326];
                
                r_data[24328] <= r_data[24327];
                
                r_data[24329] <= r_data[24328];
                
                r_data[24330] <= r_data[24329];
                
                r_data[24331] <= r_data[24330];
                
                r_data[24332] <= r_data[24331];
                
                r_data[24333] <= r_data[24332];
                
                r_data[24334] <= r_data[24333];
                
                r_data[24335] <= r_data[24334];
                
                r_data[24336] <= r_data[24335];
                
                r_data[24337] <= r_data[24336];
                
                r_data[24338] <= r_data[24337];
                
                r_data[24339] <= r_data[24338];
                
                r_data[24340] <= r_data[24339];
                
                r_data[24341] <= r_data[24340];
                
                r_data[24342] <= r_data[24341];
                
                r_data[24343] <= r_data[24342];
                
                r_data[24344] <= r_data[24343];
                
                r_data[24345] <= r_data[24344];
                
                r_data[24346] <= r_data[24345];
                
                r_data[24347] <= r_data[24346];
                
                r_data[24348] <= r_data[24347];
                
                r_data[24349] <= r_data[24348];
                
                r_data[24350] <= r_data[24349];
                
                r_data[24351] <= r_data[24350];
                
                r_data[24352] <= r_data[24351];
                
                r_data[24353] <= r_data[24352];
                
                r_data[24354] <= r_data[24353];
                
                r_data[24355] <= r_data[24354];
                
                r_data[24356] <= r_data[24355];
                
                r_data[24357] <= r_data[24356];
                
                r_data[24358] <= r_data[24357];
                
                r_data[24359] <= r_data[24358];
                
                r_data[24360] <= r_data[24359];
                
                r_data[24361] <= r_data[24360];
                
                r_data[24362] <= r_data[24361];
                
                r_data[24363] <= r_data[24362];
                
                r_data[24364] <= r_data[24363];
                
                r_data[24365] <= r_data[24364];
                
                r_data[24366] <= r_data[24365];
                
                r_data[24367] <= r_data[24366];
                
                r_data[24368] <= r_data[24367];
                
                r_data[24369] <= r_data[24368];
                
                r_data[24370] <= r_data[24369];
                
                r_data[24371] <= r_data[24370];
                
                r_data[24372] <= r_data[24371];
                
                r_data[24373] <= r_data[24372];
                
                r_data[24374] <= r_data[24373];
                
                r_data[24375] <= r_data[24374];
                
                r_data[24376] <= r_data[24375];
                
                r_data[24377] <= r_data[24376];
                
                r_data[24378] <= r_data[24377];
                
                r_data[24379] <= r_data[24378];
                
                r_data[24380] <= r_data[24379];
                
                r_data[24381] <= r_data[24380];
                
                r_data[24382] <= r_data[24381];
                
                r_data[24383] <= r_data[24382];
                
                r_data[24384] <= r_data[24383];
                
                r_data[24385] <= r_data[24384];
                
                r_data[24386] <= r_data[24385];
                
                r_data[24387] <= r_data[24386];
                
                r_data[24388] <= r_data[24387];
                
                r_data[24389] <= r_data[24388];
                
                r_data[24390] <= r_data[24389];
                
                r_data[24391] <= r_data[24390];
                
                r_data[24392] <= r_data[24391];
                
                r_data[24393] <= r_data[24392];
                
                r_data[24394] <= r_data[24393];
                
                r_data[24395] <= r_data[24394];
                
                r_data[24396] <= r_data[24395];
                
                r_data[24397] <= r_data[24396];
                
                r_data[24398] <= r_data[24397];
                
                r_data[24399] <= r_data[24398];
                
                r_data[24400] <= r_data[24399];
                
                r_data[24401] <= r_data[24400];
                
                r_data[24402] <= r_data[24401];
                
                r_data[24403] <= r_data[24402];
                
                r_data[24404] <= r_data[24403];
                
                r_data[24405] <= r_data[24404];
                
                r_data[24406] <= r_data[24405];
                
                r_data[24407] <= r_data[24406];
                
                r_data[24408] <= r_data[24407];
                
                r_data[24409] <= r_data[24408];
                
                r_data[24410] <= r_data[24409];
                
                r_data[24411] <= r_data[24410];
                
                r_data[24412] <= r_data[24411];
                
                r_data[24413] <= r_data[24412];
                
                r_data[24414] <= r_data[24413];
                
                r_data[24415] <= r_data[24414];
                
                r_data[24416] <= r_data[24415];
                
                r_data[24417] <= r_data[24416];
                
                r_data[24418] <= r_data[24417];
                
                r_data[24419] <= r_data[24418];
                
                r_data[24420] <= r_data[24419];
                
                r_data[24421] <= r_data[24420];
                
                r_data[24422] <= r_data[24421];
                
                r_data[24423] <= r_data[24422];
                
                r_data[24424] <= r_data[24423];
                
                r_data[24425] <= r_data[24424];
                
                r_data[24426] <= r_data[24425];
                
                r_data[24427] <= r_data[24426];
                
                r_data[24428] <= r_data[24427];
                
                r_data[24429] <= r_data[24428];
                
                r_data[24430] <= r_data[24429];
                
                r_data[24431] <= r_data[24430];
                
                r_data[24432] <= r_data[24431];
                
                r_data[24433] <= r_data[24432];
                
                r_data[24434] <= r_data[24433];
                
                r_data[24435] <= r_data[24434];
                
                r_data[24436] <= r_data[24435];
                
                r_data[24437] <= r_data[24436];
                
                r_data[24438] <= r_data[24437];
                
                r_data[24439] <= r_data[24438];
                
                r_data[24440] <= r_data[24439];
                
                r_data[24441] <= r_data[24440];
                
                r_data[24442] <= r_data[24441];
                
                r_data[24443] <= r_data[24442];
                
                r_data[24444] <= r_data[24443];
                
                r_data[24445] <= r_data[24444];
                
                r_data[24446] <= r_data[24445];
                
                r_data[24447] <= r_data[24446];
                
                r_data[24448] <= r_data[24447];
                
                r_data[24449] <= r_data[24448];
                
                r_data[24450] <= r_data[24449];
                
                r_data[24451] <= r_data[24450];
                
                r_data[24452] <= r_data[24451];
                
                r_data[24453] <= r_data[24452];
                
                r_data[24454] <= r_data[24453];
                
                r_data[24455] <= r_data[24454];
                
                r_data[24456] <= r_data[24455];
                
                r_data[24457] <= r_data[24456];
                
                r_data[24458] <= r_data[24457];
                
                r_data[24459] <= r_data[24458];
                
                r_data[24460] <= r_data[24459];
                
                r_data[24461] <= r_data[24460];
                
                r_data[24462] <= r_data[24461];
                
                r_data[24463] <= r_data[24462];
                
                r_data[24464] <= r_data[24463];
                
                r_data[24465] <= r_data[24464];
                
                r_data[24466] <= r_data[24465];
                
                r_data[24467] <= r_data[24466];
                
                r_data[24468] <= r_data[24467];
                
                r_data[24469] <= r_data[24468];
                
                r_data[24470] <= r_data[24469];
                
                r_data[24471] <= r_data[24470];
                
                r_data[24472] <= r_data[24471];
                
                r_data[24473] <= r_data[24472];
                
                r_data[24474] <= r_data[24473];
                
                r_data[24475] <= r_data[24474];
                
                r_data[24476] <= r_data[24475];
                
                r_data[24477] <= r_data[24476];
                
                r_data[24478] <= r_data[24477];
                
                r_data[24479] <= r_data[24478];
                
                r_data[24480] <= r_data[24479];
                
                r_data[24481] <= r_data[24480];
                
                r_data[24482] <= r_data[24481];
                
                r_data[24483] <= r_data[24482];
                
                r_data[24484] <= r_data[24483];
                
                r_data[24485] <= r_data[24484];
                
                r_data[24486] <= r_data[24485];
                
                r_data[24487] <= r_data[24486];
                
                r_data[24488] <= r_data[24487];
                
                r_data[24489] <= r_data[24488];
                
                r_data[24490] <= r_data[24489];
                
                r_data[24491] <= r_data[24490];
                
                r_data[24492] <= r_data[24491];
                
                r_data[24493] <= r_data[24492];
                
                r_data[24494] <= r_data[24493];
                
                r_data[24495] <= r_data[24494];
                
                r_data[24496] <= r_data[24495];
                
                r_data[24497] <= r_data[24496];
                
                r_data[24498] <= r_data[24497];
                
                r_data[24499] <= r_data[24498];
                
                r_data[24500] <= r_data[24499];
                
                r_data[24501] <= r_data[24500];
                
                r_data[24502] <= r_data[24501];
                
                r_data[24503] <= r_data[24502];
                
                r_data[24504] <= r_data[24503];
                
                r_data[24505] <= r_data[24504];
                
                r_data[24506] <= r_data[24505];
                
                r_data[24507] <= r_data[24506];
                
                r_data[24508] <= r_data[24507];
                
                r_data[24509] <= r_data[24508];
                
                r_data[24510] <= r_data[24509];
                
                r_data[24511] <= r_data[24510];
                
                r_data[24512] <= r_data[24511];
                
                r_data[24513] <= r_data[24512];
                
                r_data[24514] <= r_data[24513];
                
                r_data[24515] <= r_data[24514];
                
                r_data[24516] <= r_data[24515];
                
                r_data[24517] <= r_data[24516];
                
                r_data[24518] <= r_data[24517];
                
                r_data[24519] <= r_data[24518];
                
                r_data[24520] <= r_data[24519];
                
                r_data[24521] <= r_data[24520];
                
                r_data[24522] <= r_data[24521];
                
                r_data[24523] <= r_data[24522];
                
                r_data[24524] <= r_data[24523];
                
                r_data[24525] <= r_data[24524];
                
                r_data[24526] <= r_data[24525];
                
                r_data[24527] <= r_data[24526];
                
                r_data[24528] <= r_data[24527];
                
                r_data[24529] <= r_data[24528];
                
                r_data[24530] <= r_data[24529];
                
                r_data[24531] <= r_data[24530];
                
                r_data[24532] <= r_data[24531];
                
                r_data[24533] <= r_data[24532];
                
                r_data[24534] <= r_data[24533];
                
                r_data[24535] <= r_data[24534];
                
                r_data[24536] <= r_data[24535];
                
                r_data[24537] <= r_data[24536];
                
                r_data[24538] <= r_data[24537];
                
                r_data[24539] <= r_data[24538];
                
                r_data[24540] <= r_data[24539];
                
                r_data[24541] <= r_data[24540];
                
                r_data[24542] <= r_data[24541];
                
                r_data[24543] <= r_data[24542];
                
                r_data[24544] <= r_data[24543];
                
                r_data[24545] <= r_data[24544];
                
                r_data[24546] <= r_data[24545];
                
                r_data[24547] <= r_data[24546];
                
                r_data[24548] <= r_data[24547];
                
                r_data[24549] <= r_data[24548];
                
                r_data[24550] <= r_data[24549];
                
                r_data[24551] <= r_data[24550];
                
                r_data[24552] <= r_data[24551];
                
                r_data[24553] <= r_data[24552];
                
                r_data[24554] <= r_data[24553];
                
                r_data[24555] <= r_data[24554];
                
                r_data[24556] <= r_data[24555];
                
                r_data[24557] <= r_data[24556];
                
                r_data[24558] <= r_data[24557];
                
                r_data[24559] <= r_data[24558];
                
                r_data[24560] <= r_data[24559];
                
                r_data[24561] <= r_data[24560];
                
                r_data[24562] <= r_data[24561];
                
                r_data[24563] <= r_data[24562];
                
                r_data[24564] <= r_data[24563];
                
                r_data[24565] <= r_data[24564];
                
                r_data[24566] <= r_data[24565];
                
                r_data[24567] <= r_data[24566];
                
                r_data[24568] <= r_data[24567];
                
                r_data[24569] <= r_data[24568];
                
                r_data[24570] <= r_data[24569];
                
                r_data[24571] <= r_data[24570];
                
                r_data[24572] <= r_data[24571];
                
                r_data[24573] <= r_data[24572];
                
                r_data[24574] <= r_data[24573];
                
                r_data[24575] <= r_data[24574];
                
                r_data[24576] <= r_data[24575];
                
                r_data[24577] <= r_data[24576];
                
                r_data[24578] <= r_data[24577];
                
                r_data[24579] <= r_data[24578];
                
                r_data[24580] <= r_data[24579];
                
                r_data[24581] <= r_data[24580];
                
                r_data[24582] <= r_data[24581];
                
                r_data[24583] <= r_data[24582];
                
                r_data[24584] <= r_data[24583];
                
                r_data[24585] <= r_data[24584];
                
                r_data[24586] <= r_data[24585];
                
                r_data[24587] <= r_data[24586];
                
                r_data[24588] <= r_data[24587];
                
                r_data[24589] <= r_data[24588];
                
                r_data[24590] <= r_data[24589];
                
                r_data[24591] <= r_data[24590];
                
                r_data[24592] <= r_data[24591];
                
                r_data[24593] <= r_data[24592];
                
                r_data[24594] <= r_data[24593];
                
                r_data[24595] <= r_data[24594];
                
                r_data[24596] <= r_data[24595];
                
                r_data[24597] <= r_data[24596];
                
                r_data[24598] <= r_data[24597];
                
                r_data[24599] <= r_data[24598];
                
                r_data[24600] <= r_data[24599];
                
                r_data[24601] <= r_data[24600];
                
                r_data[24602] <= r_data[24601];
                
                r_data[24603] <= r_data[24602];
                
                r_data[24604] <= r_data[24603];
                
                r_data[24605] <= r_data[24604];
                
                r_data[24606] <= r_data[24605];
                
                r_data[24607] <= r_data[24606];
                
                r_data[24608] <= r_data[24607];
                
                r_data[24609] <= r_data[24608];
                
                r_data[24610] <= r_data[24609];
                
                r_data[24611] <= r_data[24610];
                
                r_data[24612] <= r_data[24611];
                
                r_data[24613] <= r_data[24612];
                
                r_data[24614] <= r_data[24613];
                
                r_data[24615] <= r_data[24614];
                
                r_data[24616] <= r_data[24615];
                
                r_data[24617] <= r_data[24616];
                
                r_data[24618] <= r_data[24617];
                
                r_data[24619] <= r_data[24618];
                
                r_data[24620] <= r_data[24619];
                
                r_data[24621] <= r_data[24620];
                
                r_data[24622] <= r_data[24621];
                
                r_data[24623] <= r_data[24622];
                
                r_data[24624] <= r_data[24623];
                
                r_data[24625] <= r_data[24624];
                
                r_data[24626] <= r_data[24625];
                
                r_data[24627] <= r_data[24626];
                
                r_data[24628] <= r_data[24627];
                
                r_data[24629] <= r_data[24628];
                
                r_data[24630] <= r_data[24629];
                
                r_data[24631] <= r_data[24630];
                
                r_data[24632] <= r_data[24631];
                
                r_data[24633] <= r_data[24632];
                
                r_data[24634] <= r_data[24633];
                
                r_data[24635] <= r_data[24634];
                
                r_data[24636] <= r_data[24635];
                
                r_data[24637] <= r_data[24636];
                
                r_data[24638] <= r_data[24637];
                
                r_data[24639] <= r_data[24638];
                
                r_data[24640] <= r_data[24639];
                
                r_data[24641] <= r_data[24640];
                
                r_data[24642] <= r_data[24641];
                
                r_data[24643] <= r_data[24642];
                
                r_data[24644] <= r_data[24643];
                
                r_data[24645] <= r_data[24644];
                
                r_data[24646] <= r_data[24645];
                
                r_data[24647] <= r_data[24646];
                
                r_data[24648] <= r_data[24647];
                
                r_data[24649] <= r_data[24648];
                
                r_data[24650] <= r_data[24649];
                
                r_data[24651] <= r_data[24650];
                
                r_data[24652] <= r_data[24651];
                
                r_data[24653] <= r_data[24652];
                
                r_data[24654] <= r_data[24653];
                
                r_data[24655] <= r_data[24654];
                
                r_data[24656] <= r_data[24655];
                
                r_data[24657] <= r_data[24656];
                
                r_data[24658] <= r_data[24657];
                
                r_data[24659] <= r_data[24658];
                
                r_data[24660] <= r_data[24659];
                
                r_data[24661] <= r_data[24660];
                
                r_data[24662] <= r_data[24661];
                
                r_data[24663] <= r_data[24662];
                
                r_data[24664] <= r_data[24663];
                
                r_data[24665] <= r_data[24664];
                
                r_data[24666] <= r_data[24665];
                
                r_data[24667] <= r_data[24666];
                
                r_data[24668] <= r_data[24667];
                
                r_data[24669] <= r_data[24668];
                
                r_data[24670] <= r_data[24669];
                
                r_data[24671] <= r_data[24670];
                
                r_data[24672] <= r_data[24671];
                
                r_data[24673] <= r_data[24672];
                
                r_data[24674] <= r_data[24673];
                
                r_data[24675] <= r_data[24674];
                
                r_data[24676] <= r_data[24675];
                
                r_data[24677] <= r_data[24676];
                
                r_data[24678] <= r_data[24677];
                
                r_data[24679] <= r_data[24678];
                
                r_data[24680] <= r_data[24679];
                
                r_data[24681] <= r_data[24680];
                
                r_data[24682] <= r_data[24681];
                
                r_data[24683] <= r_data[24682];
                
                r_data[24684] <= r_data[24683];
                
                r_data[24685] <= r_data[24684];
                
                r_data[24686] <= r_data[24685];
                
                r_data[24687] <= r_data[24686];
                
                r_data[24688] <= r_data[24687];
                
                r_data[24689] <= r_data[24688];
                
                r_data[24690] <= r_data[24689];
                
                r_data[24691] <= r_data[24690];
                
                r_data[24692] <= r_data[24691];
                
                r_data[24693] <= r_data[24692];
                
                r_data[24694] <= r_data[24693];
                
                r_data[24695] <= r_data[24694];
                
                r_data[24696] <= r_data[24695];
                
                r_data[24697] <= r_data[24696];
                
                r_data[24698] <= r_data[24697];
                
                r_data[24699] <= r_data[24698];
                
                r_data[24700] <= r_data[24699];
                
                r_data[24701] <= r_data[24700];
                
                r_data[24702] <= r_data[24701];
                
                r_data[24703] <= r_data[24702];
                
                r_data[24704] <= r_data[24703];
                
                r_data[24705] <= r_data[24704];
                
                r_data[24706] <= r_data[24705];
                
                r_data[24707] <= r_data[24706];
                
                r_data[24708] <= r_data[24707];
                
                r_data[24709] <= r_data[24708];
                
                r_data[24710] <= r_data[24709];
                
                r_data[24711] <= r_data[24710];
                
                r_data[24712] <= r_data[24711];
                
                r_data[24713] <= r_data[24712];
                
                r_data[24714] <= r_data[24713];
                
                r_data[24715] <= r_data[24714];
                
                r_data[24716] <= r_data[24715];
                
                r_data[24717] <= r_data[24716];
                
                r_data[24718] <= r_data[24717];
                
                r_data[24719] <= r_data[24718];
                
                r_data[24720] <= r_data[24719];
                
                r_data[24721] <= r_data[24720];
                
                r_data[24722] <= r_data[24721];
                
                r_data[24723] <= r_data[24722];
                
                r_data[24724] <= r_data[24723];
                
                r_data[24725] <= r_data[24724];
                
                r_data[24726] <= r_data[24725];
                
                r_data[24727] <= r_data[24726];
                
                r_data[24728] <= r_data[24727];
                
                r_data[24729] <= r_data[24728];
                
                r_data[24730] <= r_data[24729];
                
                r_data[24731] <= r_data[24730];
                
                r_data[24732] <= r_data[24731];
                
                r_data[24733] <= r_data[24732];
                
                r_data[24734] <= r_data[24733];
                
                r_data[24735] <= r_data[24734];
                
                r_data[24736] <= r_data[24735];
                
                r_data[24737] <= r_data[24736];
                
                r_data[24738] <= r_data[24737];
                
                r_data[24739] <= r_data[24738];
                
                r_data[24740] <= r_data[24739];
                
                r_data[24741] <= r_data[24740];
                
                r_data[24742] <= r_data[24741];
                
                r_data[24743] <= r_data[24742];
                
                r_data[24744] <= r_data[24743];
                
                r_data[24745] <= r_data[24744];
                
                r_data[24746] <= r_data[24745];
                
                r_data[24747] <= r_data[24746];
                
                r_data[24748] <= r_data[24747];
                
                r_data[24749] <= r_data[24748];
                
                r_data[24750] <= r_data[24749];
                
                r_data[24751] <= r_data[24750];
                
                r_data[24752] <= r_data[24751];
                
                r_data[24753] <= r_data[24752];
                
                r_data[24754] <= r_data[24753];
                
                r_data[24755] <= r_data[24754];
                
                r_data[24756] <= r_data[24755];
                
                r_data[24757] <= r_data[24756];
                
                r_data[24758] <= r_data[24757];
                
                r_data[24759] <= r_data[24758];
                
                r_data[24760] <= r_data[24759];
                
                r_data[24761] <= r_data[24760];
                
                r_data[24762] <= r_data[24761];
                
                r_data[24763] <= r_data[24762];
                
                r_data[24764] <= r_data[24763];
                
                r_data[24765] <= r_data[24764];
                
                r_data[24766] <= r_data[24765];
                
                r_data[24767] <= r_data[24766];
                
                r_data[24768] <= r_data[24767];
                
                r_data[24769] <= r_data[24768];
                
                r_data[24770] <= r_data[24769];
                
                r_data[24771] <= r_data[24770];
                
                r_data[24772] <= r_data[24771];
                
                r_data[24773] <= r_data[24772];
                
                r_data[24774] <= r_data[24773];
                
                r_data[24775] <= r_data[24774];
                
                r_data[24776] <= r_data[24775];
                
                r_data[24777] <= r_data[24776];
                
                r_data[24778] <= r_data[24777];
                
                r_data[24779] <= r_data[24778];
                
                r_data[24780] <= r_data[24779];
                
                r_data[24781] <= r_data[24780];
                
                r_data[24782] <= r_data[24781];
                
                r_data[24783] <= r_data[24782];
                
                r_data[24784] <= r_data[24783];
                
                r_data[24785] <= r_data[24784];
                
                r_data[24786] <= r_data[24785];
                
                r_data[24787] <= r_data[24786];
                
                r_data[24788] <= r_data[24787];
                
                r_data[24789] <= r_data[24788];
                
                r_data[24790] <= r_data[24789];
                
                r_data[24791] <= r_data[24790];
                
                r_data[24792] <= r_data[24791];
                
                r_data[24793] <= r_data[24792];
                
                r_data[24794] <= r_data[24793];
                
                r_data[24795] <= r_data[24794];
                
                r_data[24796] <= r_data[24795];
                
                r_data[24797] <= r_data[24796];
                
                r_data[24798] <= r_data[24797];
                
                r_data[24799] <= r_data[24798];
                
                r_data[24800] <= r_data[24799];
                
                r_data[24801] <= r_data[24800];
                
                r_data[24802] <= r_data[24801];
                
                r_data[24803] <= r_data[24802];
                
                r_data[24804] <= r_data[24803];
                
                r_data[24805] <= r_data[24804];
                
                r_data[24806] <= r_data[24805];
                
                r_data[24807] <= r_data[24806];
                
                r_data[24808] <= r_data[24807];
                
                r_data[24809] <= r_data[24808];
                
                r_data[24810] <= r_data[24809];
                
                r_data[24811] <= r_data[24810];
                
                r_data[24812] <= r_data[24811];
                
                r_data[24813] <= r_data[24812];
                
                r_data[24814] <= r_data[24813];
                
                r_data[24815] <= r_data[24814];
                
                r_data[24816] <= r_data[24815];
                
                r_data[24817] <= r_data[24816];
                
                r_data[24818] <= r_data[24817];
                
                r_data[24819] <= r_data[24818];
                
                r_data[24820] <= r_data[24819];
                
                r_data[24821] <= r_data[24820];
                
                r_data[24822] <= r_data[24821];
                
                r_data[24823] <= r_data[24822];
                
                r_data[24824] <= r_data[24823];
                
                r_data[24825] <= r_data[24824];
                
                r_data[24826] <= r_data[24825];
                
                r_data[24827] <= r_data[24826];
                
                r_data[24828] <= r_data[24827];
                
                r_data[24829] <= r_data[24828];
                
                r_data[24830] <= r_data[24829];
                
                r_data[24831] <= r_data[24830];
                
                r_data[24832] <= r_data[24831];
                
                r_data[24833] <= r_data[24832];
                
                r_data[24834] <= r_data[24833];
                
                r_data[24835] <= r_data[24834];
                
                r_data[24836] <= r_data[24835];
                
                r_data[24837] <= r_data[24836];
                
                r_data[24838] <= r_data[24837];
                
                r_data[24839] <= r_data[24838];
                
                r_data[24840] <= r_data[24839];
                
                r_data[24841] <= r_data[24840];
                
                r_data[24842] <= r_data[24841];
                
                r_data[24843] <= r_data[24842];
                
                r_data[24844] <= r_data[24843];
                
                r_data[24845] <= r_data[24844];
                
                r_data[24846] <= r_data[24845];
                
                r_data[24847] <= r_data[24846];
                
                r_data[24848] <= r_data[24847];
                
                r_data[24849] <= r_data[24848];
                
                r_data[24850] <= r_data[24849];
                
                r_data[24851] <= r_data[24850];
                
                r_data[24852] <= r_data[24851];
                
                r_data[24853] <= r_data[24852];
                
                r_data[24854] <= r_data[24853];
                
                r_data[24855] <= r_data[24854];
                
                r_data[24856] <= r_data[24855];
                
                r_data[24857] <= r_data[24856];
                
                r_data[24858] <= r_data[24857];
                
                r_data[24859] <= r_data[24858];
                
                r_data[24860] <= r_data[24859];
                
                r_data[24861] <= r_data[24860];
                
                r_data[24862] <= r_data[24861];
                
                r_data[24863] <= r_data[24862];
                
                r_data[24864] <= r_data[24863];
                
                r_data[24865] <= r_data[24864];
                
                r_data[24866] <= r_data[24865];
                
                r_data[24867] <= r_data[24866];
                
                r_data[24868] <= r_data[24867];
                
                r_data[24869] <= r_data[24868];
                
                r_data[24870] <= r_data[24869];
                
                r_data[24871] <= r_data[24870];
                
                r_data[24872] <= r_data[24871];
                
                r_data[24873] <= r_data[24872];
                
                r_data[24874] <= r_data[24873];
                
                r_data[24875] <= r_data[24874];
                
                r_data[24876] <= r_data[24875];
                
                r_data[24877] <= r_data[24876];
                
                r_data[24878] <= r_data[24877];
                
                r_data[24879] <= r_data[24878];
                
                r_data[24880] <= r_data[24879];
                
                r_data[24881] <= r_data[24880];
                
                r_data[24882] <= r_data[24881];
                
                r_data[24883] <= r_data[24882];
                
                r_data[24884] <= r_data[24883];
                
                r_data[24885] <= r_data[24884];
                
                r_data[24886] <= r_data[24885];
                
                r_data[24887] <= r_data[24886];
                
                r_data[24888] <= r_data[24887];
                
                r_data[24889] <= r_data[24888];
                
                r_data[24890] <= r_data[24889];
                
                r_data[24891] <= r_data[24890];
                
                r_data[24892] <= r_data[24891];
                
                r_data[24893] <= r_data[24892];
                
                r_data[24894] <= r_data[24893];
                
                r_data[24895] <= r_data[24894];
                
                r_data[24896] <= r_data[24895];
                
                r_data[24897] <= r_data[24896];
                
                r_data[24898] <= r_data[24897];
                
                r_data[24899] <= r_data[24898];
                
                r_data[24900] <= r_data[24899];
                
                r_data[24901] <= r_data[24900];
                
                r_data[24902] <= r_data[24901];
                
                r_data[24903] <= r_data[24902];
                
                r_data[24904] <= r_data[24903];
                
                r_data[24905] <= r_data[24904];
                
                r_data[24906] <= r_data[24905];
                
                r_data[24907] <= r_data[24906];
                
                r_data[24908] <= r_data[24907];
                
                r_data[24909] <= r_data[24908];
                
                r_data[24910] <= r_data[24909];
                
                r_data[24911] <= r_data[24910];
                
                r_data[24912] <= r_data[24911];
                
                r_data[24913] <= r_data[24912];
                
                r_data[24914] <= r_data[24913];
                
                r_data[24915] <= r_data[24914];
                
                r_data[24916] <= r_data[24915];
                
                r_data[24917] <= r_data[24916];
                
                r_data[24918] <= r_data[24917];
                
                r_data[24919] <= r_data[24918];
                
                r_data[24920] <= r_data[24919];
                
                r_data[24921] <= r_data[24920];
                
                r_data[24922] <= r_data[24921];
                
                r_data[24923] <= r_data[24922];
                
                r_data[24924] <= r_data[24923];
                
                r_data[24925] <= r_data[24924];
                
                r_data[24926] <= r_data[24925];
                
                r_data[24927] <= r_data[24926];
                
                r_data[24928] <= r_data[24927];
                
                r_data[24929] <= r_data[24928];
                
                r_data[24930] <= r_data[24929];
                
                r_data[24931] <= r_data[24930];
                
                r_data[24932] <= r_data[24931];
                
                r_data[24933] <= r_data[24932];
                
                r_data[24934] <= r_data[24933];
                
                r_data[24935] <= r_data[24934];
                
                r_data[24936] <= r_data[24935];
                
                r_data[24937] <= r_data[24936];
                
                r_data[24938] <= r_data[24937];
                
                r_data[24939] <= r_data[24938];
                
                r_data[24940] <= r_data[24939];
                
                r_data[24941] <= r_data[24940];
                
                r_data[24942] <= r_data[24941];
                
                r_data[24943] <= r_data[24942];
                
                r_data[24944] <= r_data[24943];
                
                r_data[24945] <= r_data[24944];
                
                r_data[24946] <= r_data[24945];
                
                r_data[24947] <= r_data[24946];
                
                r_data[24948] <= r_data[24947];
                
                r_data[24949] <= r_data[24948];
                
                r_data[24950] <= r_data[24949];
                
                r_data[24951] <= r_data[24950];
                
                r_data[24952] <= r_data[24951];
                
                r_data[24953] <= r_data[24952];
                
                r_data[24954] <= r_data[24953];
                
                r_data[24955] <= r_data[24954];
                
                r_data[24956] <= r_data[24955];
                
                r_data[24957] <= r_data[24956];
                
                r_data[24958] <= r_data[24957];
                
                r_data[24959] <= r_data[24958];
                
                r_data[24960] <= r_data[24959];
                
                r_data[24961] <= r_data[24960];
                
                r_data[24962] <= r_data[24961];
                
                r_data[24963] <= r_data[24962];
                
                r_data[24964] <= r_data[24963];
                
                r_data[24965] <= r_data[24964];
                
                r_data[24966] <= r_data[24965];
                
                r_data[24967] <= r_data[24966];
                
                r_data[24968] <= r_data[24967];
                
                r_data[24969] <= r_data[24968];
                
                r_data[24970] <= r_data[24969];
                
                r_data[24971] <= r_data[24970];
                
                r_data[24972] <= r_data[24971];
                
                r_data[24973] <= r_data[24972];
                
                r_data[24974] <= r_data[24973];
                
                r_data[24975] <= r_data[24974];
                
                r_data[24976] <= r_data[24975];
                
                r_data[24977] <= r_data[24976];
                
                r_data[24978] <= r_data[24977];
                
                r_data[24979] <= r_data[24978];
                
                r_data[24980] <= r_data[24979];
                
                r_data[24981] <= r_data[24980];
                
                r_data[24982] <= r_data[24981];
                
                r_data[24983] <= r_data[24982];
                
                r_data[24984] <= r_data[24983];
                
                r_data[24985] <= r_data[24984];
                
                r_data[24986] <= r_data[24985];
                
                r_data[24987] <= r_data[24986];
                
                r_data[24988] <= r_data[24987];
                
                r_data[24989] <= r_data[24988];
                
                r_data[24990] <= r_data[24989];
                
                r_data[24991] <= r_data[24990];
                
                r_data[24992] <= r_data[24991];
                
                r_data[24993] <= r_data[24992];
                
                r_data[24994] <= r_data[24993];
                
                r_data[24995] <= r_data[24994];
                
                r_data[24996] <= r_data[24995];
                
                r_data[24997] <= r_data[24996];
                
                r_data[24998] <= r_data[24997];
                
                r_data[24999] <= r_data[24998];
                
                r_data[25000] <= r_data[24999];
                
                r_data[25001] <= r_data[25000];
                
                r_data[25002] <= r_data[25001];
                
                r_data[25003] <= r_data[25002];
                
                r_data[25004] <= r_data[25003];
                
                r_data[25005] <= r_data[25004];
                
                r_data[25006] <= r_data[25005];
                
                r_data[25007] <= r_data[25006];
                
                r_data[25008] <= r_data[25007];
                
                r_data[25009] <= r_data[25008];
                
                r_data[25010] <= r_data[25009];
                
                r_data[25011] <= r_data[25010];
                
                r_data[25012] <= r_data[25011];
                
                r_data[25013] <= r_data[25012];
                
                r_data[25014] <= r_data[25013];
                
                r_data[25015] <= r_data[25014];
                
                r_data[25016] <= r_data[25015];
                
                r_data[25017] <= r_data[25016];
                
                r_data[25018] <= r_data[25017];
                
                r_data[25019] <= r_data[25018];
                
                r_data[25020] <= r_data[25019];
                
                r_data[25021] <= r_data[25020];
                
                r_data[25022] <= r_data[25021];
                
                r_data[25023] <= r_data[25022];
                
                r_data[25024] <= r_data[25023];
                
                r_data[25025] <= r_data[25024];
                
                r_data[25026] <= r_data[25025];
                
                r_data[25027] <= r_data[25026];
                
                r_data[25028] <= r_data[25027];
                
                r_data[25029] <= r_data[25028];
                
                r_data[25030] <= r_data[25029];
                
                r_data[25031] <= r_data[25030];
                
                r_data[25032] <= r_data[25031];
                
                r_data[25033] <= r_data[25032];
                
                r_data[25034] <= r_data[25033];
                
                r_data[25035] <= r_data[25034];
                
                r_data[25036] <= r_data[25035];
                
                r_data[25037] <= r_data[25036];
                
                r_data[25038] <= r_data[25037];
                
                r_data[25039] <= r_data[25038];
                
                r_data[25040] <= r_data[25039];
                
                r_data[25041] <= r_data[25040];
                
                r_data[25042] <= r_data[25041];
                
                r_data[25043] <= r_data[25042];
                
                r_data[25044] <= r_data[25043];
                
                r_data[25045] <= r_data[25044];
                
                r_data[25046] <= r_data[25045];
                
                r_data[25047] <= r_data[25046];
                
                r_data[25048] <= r_data[25047];
                
                r_data[25049] <= r_data[25048];
                
                r_data[25050] <= r_data[25049];
                
                r_data[25051] <= r_data[25050];
                
                r_data[25052] <= r_data[25051];
                
                r_data[25053] <= r_data[25052];
                
                r_data[25054] <= r_data[25053];
                
                r_data[25055] <= r_data[25054];
                
                r_data[25056] <= r_data[25055];
                
                r_data[25057] <= r_data[25056];
                
                r_data[25058] <= r_data[25057];
                
                r_data[25059] <= r_data[25058];
                
                r_data[25060] <= r_data[25059];
                
                r_data[25061] <= r_data[25060];
                
                r_data[25062] <= r_data[25061];
                
                r_data[25063] <= r_data[25062];
                
                r_data[25064] <= r_data[25063];
                
                r_data[25065] <= r_data[25064];
                
                r_data[25066] <= r_data[25065];
                
                r_data[25067] <= r_data[25066];
                
                r_data[25068] <= r_data[25067];
                
                r_data[25069] <= r_data[25068];
                
                r_data[25070] <= r_data[25069];
                
                r_data[25071] <= r_data[25070];
                
                r_data[25072] <= r_data[25071];
                
                r_data[25073] <= r_data[25072];
                
                r_data[25074] <= r_data[25073];
                
                r_data[25075] <= r_data[25074];
                
                r_data[25076] <= r_data[25075];
                
                r_data[25077] <= r_data[25076];
                
                r_data[25078] <= r_data[25077];
                
                r_data[25079] <= r_data[25078];
                
                r_data[25080] <= r_data[25079];
                
                r_data[25081] <= r_data[25080];
                
                r_data[25082] <= r_data[25081];
                
                r_data[25083] <= r_data[25082];
                
                r_data[25084] <= r_data[25083];
                
                r_data[25085] <= r_data[25084];
                
                r_data[25086] <= r_data[25085];
                
                r_data[25087] <= r_data[25086];
                
                r_data[25088] <= r_data[25087];
                
                r_data[25089] <= r_data[25088];
                
                r_data[25090] <= r_data[25089];
                
                r_data[25091] <= r_data[25090];
                
                r_data[25092] <= r_data[25091];
                
                r_data[25093] <= r_data[25092];
                
                r_data[25094] <= r_data[25093];
                
                r_data[25095] <= r_data[25094];
                
                r_data[25096] <= r_data[25095];
                
                r_data[25097] <= r_data[25096];
                
                r_data[25098] <= r_data[25097];
                
                r_data[25099] <= r_data[25098];
                
                r_data[25100] <= r_data[25099];
                
                r_data[25101] <= r_data[25100];
                
                r_data[25102] <= r_data[25101];
                
                r_data[25103] <= r_data[25102];
                
                r_data[25104] <= r_data[25103];
                
                r_data[25105] <= r_data[25104];
                
                r_data[25106] <= r_data[25105];
                
                r_data[25107] <= r_data[25106];
                
                r_data[25108] <= r_data[25107];
                
                r_data[25109] <= r_data[25108];
                
                r_data[25110] <= r_data[25109];
                
                r_data[25111] <= r_data[25110];
                
                r_data[25112] <= r_data[25111];
                
                r_data[25113] <= r_data[25112];
                
                r_data[25114] <= r_data[25113];
                
                r_data[25115] <= r_data[25114];
                
                r_data[25116] <= r_data[25115];
                
                r_data[25117] <= r_data[25116];
                
                r_data[25118] <= r_data[25117];
                
                r_data[25119] <= r_data[25118];
                
                r_data[25120] <= r_data[25119];
                
                r_data[25121] <= r_data[25120];
                
                r_data[25122] <= r_data[25121];
                
                r_data[25123] <= r_data[25122];
                
                r_data[25124] <= r_data[25123];
                
                r_data[25125] <= r_data[25124];
                
                r_data[25126] <= r_data[25125];
                
                r_data[25127] <= r_data[25126];
                
                r_data[25128] <= r_data[25127];
                
                r_data[25129] <= r_data[25128];
                
                r_data[25130] <= r_data[25129];
                
                r_data[25131] <= r_data[25130];
                
                r_data[25132] <= r_data[25131];
                
                r_data[25133] <= r_data[25132];
                
                r_data[25134] <= r_data[25133];
                
                r_data[25135] <= r_data[25134];
                
                r_data[25136] <= r_data[25135];
                
                r_data[25137] <= r_data[25136];
                
                r_data[25138] <= r_data[25137];
                
                r_data[25139] <= r_data[25138];
                
                r_data[25140] <= r_data[25139];
                
                r_data[25141] <= r_data[25140];
                
                r_data[25142] <= r_data[25141];
                
                r_data[25143] <= r_data[25142];
                
                r_data[25144] <= r_data[25143];
                
                r_data[25145] <= r_data[25144];
                
                r_data[25146] <= r_data[25145];
                
                r_data[25147] <= r_data[25146];
                
                r_data[25148] <= r_data[25147];
                
                r_data[25149] <= r_data[25148];
                
                r_data[25150] <= r_data[25149];
                
                r_data[25151] <= r_data[25150];
                
                r_data[25152] <= r_data[25151];
                
                r_data[25153] <= r_data[25152];
                
                r_data[25154] <= r_data[25153];
                
                r_data[25155] <= r_data[25154];
                
                r_data[25156] <= r_data[25155];
                
                r_data[25157] <= r_data[25156];
                
                r_data[25158] <= r_data[25157];
                
                r_data[25159] <= r_data[25158];
                
                r_data[25160] <= r_data[25159];
                
                r_data[25161] <= r_data[25160];
                
                r_data[25162] <= r_data[25161];
                
                r_data[25163] <= r_data[25162];
                
                r_data[25164] <= r_data[25163];
                
                r_data[25165] <= r_data[25164];
                
                r_data[25166] <= r_data[25165];
                
                r_data[25167] <= r_data[25166];
                
                r_data[25168] <= r_data[25167];
                
                r_data[25169] <= r_data[25168];
                
                r_data[25170] <= r_data[25169];
                
                r_data[25171] <= r_data[25170];
                
                r_data[25172] <= r_data[25171];
                
                r_data[25173] <= r_data[25172];
                
                r_data[25174] <= r_data[25173];
                
                r_data[25175] <= r_data[25174];
                
                r_data[25176] <= r_data[25175];
                
                r_data[25177] <= r_data[25176];
                
                r_data[25178] <= r_data[25177];
                
                r_data[25179] <= r_data[25178];
                
                r_data[25180] <= r_data[25179];
                
                r_data[25181] <= r_data[25180];
                
                r_data[25182] <= r_data[25181];
                
                r_data[25183] <= r_data[25182];
                
                r_data[25184] <= r_data[25183];
                
                r_data[25185] <= r_data[25184];
                
                r_data[25186] <= r_data[25185];
                
                r_data[25187] <= r_data[25186];
                
                r_data[25188] <= r_data[25187];
                
                r_data[25189] <= r_data[25188];
                
                r_data[25190] <= r_data[25189];
                
                r_data[25191] <= r_data[25190];
                
                r_data[25192] <= r_data[25191];
                
                r_data[25193] <= r_data[25192];
                
                r_data[25194] <= r_data[25193];
                
                r_data[25195] <= r_data[25194];
                
                r_data[25196] <= r_data[25195];
                
                r_data[25197] <= r_data[25196];
                
                r_data[25198] <= r_data[25197];
                
                r_data[25199] <= r_data[25198];
                
                r_data[25200] <= r_data[25199];
                
                r_data[25201] <= r_data[25200];
                
                r_data[25202] <= r_data[25201];
                
                r_data[25203] <= r_data[25202];
                
                r_data[25204] <= r_data[25203];
                
                r_data[25205] <= r_data[25204];
                
                r_data[25206] <= r_data[25205];
                
                r_data[25207] <= r_data[25206];
                
                r_data[25208] <= r_data[25207];
                
                r_data[25209] <= r_data[25208];
                
                r_data[25210] <= r_data[25209];
                
                r_data[25211] <= r_data[25210];
                
                r_data[25212] <= r_data[25211];
                
                r_data[25213] <= r_data[25212];
                
                r_data[25214] <= r_data[25213];
                
                r_data[25215] <= r_data[25214];
                
                r_data[25216] <= r_data[25215];
                
                r_data[25217] <= r_data[25216];
                
                r_data[25218] <= r_data[25217];
                
                r_data[25219] <= r_data[25218];
                
                r_data[25220] <= r_data[25219];
                
                r_data[25221] <= r_data[25220];
                
                r_data[25222] <= r_data[25221];
                
                r_data[25223] <= r_data[25222];
                
                r_data[25224] <= r_data[25223];
                
                r_data[25225] <= r_data[25224];
                
                r_data[25226] <= r_data[25225];
                
                r_data[25227] <= r_data[25226];
                
                r_data[25228] <= r_data[25227];
                
                r_data[25229] <= r_data[25228];
                
                r_data[25230] <= r_data[25229];
                
                r_data[25231] <= r_data[25230];
                
                r_data[25232] <= r_data[25231];
                
                r_data[25233] <= r_data[25232];
                
                r_data[25234] <= r_data[25233];
                
                r_data[25235] <= r_data[25234];
                
                r_data[25236] <= r_data[25235];
                
                r_data[25237] <= r_data[25236];
                
                r_data[25238] <= r_data[25237];
                
                r_data[25239] <= r_data[25238];
                
                r_data[25240] <= r_data[25239];
                
                r_data[25241] <= r_data[25240];
                
                r_data[25242] <= r_data[25241];
                
                r_data[25243] <= r_data[25242];
                
                r_data[25244] <= r_data[25243];
                
                r_data[25245] <= r_data[25244];
                
                r_data[25246] <= r_data[25245];
                
                r_data[25247] <= r_data[25246];
                
                r_data[25248] <= r_data[25247];
                
                r_data[25249] <= r_data[25248];
                
                r_data[25250] <= r_data[25249];
                
                r_data[25251] <= r_data[25250];
                
                r_data[25252] <= r_data[25251];
                
                r_data[25253] <= r_data[25252];
                
                r_data[25254] <= r_data[25253];
                
                r_data[25255] <= r_data[25254];
                
                r_data[25256] <= r_data[25255];
                
                r_data[25257] <= r_data[25256];
                
                r_data[25258] <= r_data[25257];
                
                r_data[25259] <= r_data[25258];
                
                r_data[25260] <= r_data[25259];
                
                r_data[25261] <= r_data[25260];
                
                r_data[25262] <= r_data[25261];
                
                r_data[25263] <= r_data[25262];
                
                r_data[25264] <= r_data[25263];
                
                r_data[25265] <= r_data[25264];
                
                r_data[25266] <= r_data[25265];
                
                r_data[25267] <= r_data[25266];
                
                r_data[25268] <= r_data[25267];
                
                r_data[25269] <= r_data[25268];
                
                r_data[25270] <= r_data[25269];
                
                r_data[25271] <= r_data[25270];
                
                r_data[25272] <= r_data[25271];
                
                r_data[25273] <= r_data[25272];
                
                r_data[25274] <= r_data[25273];
                
                r_data[25275] <= r_data[25274];
                
                r_data[25276] <= r_data[25275];
                
                r_data[25277] <= r_data[25276];
                
                r_data[25278] <= r_data[25277];
                
                r_data[25279] <= r_data[25278];
                
                r_data[25280] <= r_data[25279];
                
                r_data[25281] <= r_data[25280];
                
                r_data[25282] <= r_data[25281];
                
                r_data[25283] <= r_data[25282];
                
                r_data[25284] <= r_data[25283];
                
                r_data[25285] <= r_data[25284];
                
                r_data[25286] <= r_data[25285];
                
                r_data[25287] <= r_data[25286];
                
                r_data[25288] <= r_data[25287];
                
                r_data[25289] <= r_data[25288];
                
                r_data[25290] <= r_data[25289];
                
                r_data[25291] <= r_data[25290];
                
                r_data[25292] <= r_data[25291];
                
                r_data[25293] <= r_data[25292];
                
                r_data[25294] <= r_data[25293];
                
                r_data[25295] <= r_data[25294];
                
                r_data[25296] <= r_data[25295];
                
                r_data[25297] <= r_data[25296];
                
                r_data[25298] <= r_data[25297];
                
                r_data[25299] <= r_data[25298];
                
                r_data[25300] <= r_data[25299];
                
                r_data[25301] <= r_data[25300];
                
                r_data[25302] <= r_data[25301];
                
                r_data[25303] <= r_data[25302];
                
                r_data[25304] <= r_data[25303];
                
                r_data[25305] <= r_data[25304];
                
                r_data[25306] <= r_data[25305];
                
                r_data[25307] <= r_data[25306];
                
                r_data[25308] <= r_data[25307];
                
                r_data[25309] <= r_data[25308];
                
                r_data[25310] <= r_data[25309];
                
                r_data[25311] <= r_data[25310];
                
                r_data[25312] <= r_data[25311];
                
                r_data[25313] <= r_data[25312];
                
                r_data[25314] <= r_data[25313];
                
                r_data[25315] <= r_data[25314];
                
                r_data[25316] <= r_data[25315];
                
                r_data[25317] <= r_data[25316];
                
                r_data[25318] <= r_data[25317];
                
                r_data[25319] <= r_data[25318];
                
                r_data[25320] <= r_data[25319];
                
                r_data[25321] <= r_data[25320];
                
                r_data[25322] <= r_data[25321];
                
                r_data[25323] <= r_data[25322];
                
                r_data[25324] <= r_data[25323];
                
                r_data[25325] <= r_data[25324];
                
                r_data[25326] <= r_data[25325];
                
                r_data[25327] <= r_data[25326];
                
                r_data[25328] <= r_data[25327];
                
                r_data[25329] <= r_data[25328];
                
                r_data[25330] <= r_data[25329];
                
                r_data[25331] <= r_data[25330];
                
                r_data[25332] <= r_data[25331];
                
                r_data[25333] <= r_data[25332];
                
                r_data[25334] <= r_data[25333];
                
                r_data[25335] <= r_data[25334];
                
                r_data[25336] <= r_data[25335];
                
                r_data[25337] <= r_data[25336];
                
                r_data[25338] <= r_data[25337];
                
                r_data[25339] <= r_data[25338];
                
                r_data[25340] <= r_data[25339];
                
                r_data[25341] <= r_data[25340];
                
                r_data[25342] <= r_data[25341];
                
                r_data[25343] <= r_data[25342];
                
                r_data[25344] <= r_data[25343];
                
                r_data[25345] <= r_data[25344];
                
                r_data[25346] <= r_data[25345];
                
                r_data[25347] <= r_data[25346];
                
                r_data[25348] <= r_data[25347];
                
                r_data[25349] <= r_data[25348];
                
                r_data[25350] <= r_data[25349];
                
                r_data[25351] <= r_data[25350];
                
                r_data[25352] <= r_data[25351];
                
                r_data[25353] <= r_data[25352];
                
                r_data[25354] <= r_data[25353];
                
                r_data[25355] <= r_data[25354];
                
                r_data[25356] <= r_data[25355];
                
                r_data[25357] <= r_data[25356];
                
                r_data[25358] <= r_data[25357];
                
                r_data[25359] <= r_data[25358];
                
                r_data[25360] <= r_data[25359];
                
                r_data[25361] <= r_data[25360];
                
                r_data[25362] <= r_data[25361];
                
                r_data[25363] <= r_data[25362];
                
                r_data[25364] <= r_data[25363];
                
                r_data[25365] <= r_data[25364];
                
                r_data[25366] <= r_data[25365];
                
                r_data[25367] <= r_data[25366];
                
                r_data[25368] <= r_data[25367];
                
                r_data[25369] <= r_data[25368];
                
                r_data[25370] <= r_data[25369];
                
                r_data[25371] <= r_data[25370];
                
                r_data[25372] <= r_data[25371];
                
                r_data[25373] <= r_data[25372];
                
                r_data[25374] <= r_data[25373];
                
                r_data[25375] <= r_data[25374];
                
                r_data[25376] <= r_data[25375];
                
                r_data[25377] <= r_data[25376];
                
                r_data[25378] <= r_data[25377];
                
                r_data[25379] <= r_data[25378];
                
                r_data[25380] <= r_data[25379];
                
                r_data[25381] <= r_data[25380];
                
                r_data[25382] <= r_data[25381];
                
                r_data[25383] <= r_data[25382];
                
                r_data[25384] <= r_data[25383];
                
                r_data[25385] <= r_data[25384];
                
                r_data[25386] <= r_data[25385];
                
                r_data[25387] <= r_data[25386];
                
                r_data[25388] <= r_data[25387];
                
                r_data[25389] <= r_data[25388];
                
                r_data[25390] <= r_data[25389];
                
                r_data[25391] <= r_data[25390];
                
                r_data[25392] <= r_data[25391];
                
                r_data[25393] <= r_data[25392];
                
                r_data[25394] <= r_data[25393];
                
                r_data[25395] <= r_data[25394];
                
                r_data[25396] <= r_data[25395];
                
                r_data[25397] <= r_data[25396];
                
                r_data[25398] <= r_data[25397];
                
                r_data[25399] <= r_data[25398];
                
                r_data[25400] <= r_data[25399];
                
                r_data[25401] <= r_data[25400];
                
                r_data[25402] <= r_data[25401];
                
                r_data[25403] <= r_data[25402];
                
                r_data[25404] <= r_data[25403];
                
                r_data[25405] <= r_data[25404];
                
                r_data[25406] <= r_data[25405];
                
                r_data[25407] <= r_data[25406];
                
                r_data[25408] <= r_data[25407];
                
                r_data[25409] <= r_data[25408];
                
                r_data[25410] <= r_data[25409];
                
                r_data[25411] <= r_data[25410];
                
                r_data[25412] <= r_data[25411];
                
                r_data[25413] <= r_data[25412];
                
                r_data[25414] <= r_data[25413];
                
                r_data[25415] <= r_data[25414];
                
                r_data[25416] <= r_data[25415];
                
                r_data[25417] <= r_data[25416];
                
                r_data[25418] <= r_data[25417];
                
                r_data[25419] <= r_data[25418];
                
                r_data[25420] <= r_data[25419];
                
                r_data[25421] <= r_data[25420];
                
                r_data[25422] <= r_data[25421];
                
                r_data[25423] <= r_data[25422];
                
                r_data[25424] <= r_data[25423];
                
                r_data[25425] <= r_data[25424];
                
                r_data[25426] <= r_data[25425];
                
                r_data[25427] <= r_data[25426];
                
                r_data[25428] <= r_data[25427];
                
                r_data[25429] <= r_data[25428];
                
                r_data[25430] <= r_data[25429];
                
                r_data[25431] <= r_data[25430];
                
                r_data[25432] <= r_data[25431];
                
                r_data[25433] <= r_data[25432];
                
                r_data[25434] <= r_data[25433];
                
                r_data[25435] <= r_data[25434];
                
                r_data[25436] <= r_data[25435];
                
                r_data[25437] <= r_data[25436];
                
                r_data[25438] <= r_data[25437];
                
                r_data[25439] <= r_data[25438];
                
                r_data[25440] <= r_data[25439];
                
                r_data[25441] <= r_data[25440];
                
                r_data[25442] <= r_data[25441];
                
                r_data[25443] <= r_data[25442];
                
                r_data[25444] <= r_data[25443];
                
                r_data[25445] <= r_data[25444];
                
                r_data[25446] <= r_data[25445];
                
                r_data[25447] <= r_data[25446];
                
                r_data[25448] <= r_data[25447];
                
                r_data[25449] <= r_data[25448];
                
                r_data[25450] <= r_data[25449];
                
                r_data[25451] <= r_data[25450];
                
                r_data[25452] <= r_data[25451];
                
                r_data[25453] <= r_data[25452];
                
                r_data[25454] <= r_data[25453];
                
                r_data[25455] <= r_data[25454];
                
                r_data[25456] <= r_data[25455];
                
                r_data[25457] <= r_data[25456];
                
                r_data[25458] <= r_data[25457];
                
                r_data[25459] <= r_data[25458];
                
                r_data[25460] <= r_data[25459];
                
                r_data[25461] <= r_data[25460];
                
                r_data[25462] <= r_data[25461];
                
                r_data[25463] <= r_data[25462];
                
                r_data[25464] <= r_data[25463];
                
                r_data[25465] <= r_data[25464];
                
                r_data[25466] <= r_data[25465];
                
                r_data[25467] <= r_data[25466];
                
                r_data[25468] <= r_data[25467];
                
                r_data[25469] <= r_data[25468];
                
                r_data[25470] <= r_data[25469];
                
                r_data[25471] <= r_data[25470];
                
                r_data[25472] <= r_data[25471];
                
                r_data[25473] <= r_data[25472];
                
                r_data[25474] <= r_data[25473];
                
                r_data[25475] <= r_data[25474];
                
                r_data[25476] <= r_data[25475];
                
                r_data[25477] <= r_data[25476];
                
                r_data[25478] <= r_data[25477];
                
                r_data[25479] <= r_data[25478];
                
                r_data[25480] <= r_data[25479];
                
                r_data[25481] <= r_data[25480];
                
                r_data[25482] <= r_data[25481];
                
                r_data[25483] <= r_data[25482];
                
                r_data[25484] <= r_data[25483];
                
                r_data[25485] <= r_data[25484];
                
                r_data[25486] <= r_data[25485];
                
                r_data[25487] <= r_data[25486];
                
                r_data[25488] <= r_data[25487];
                
                r_data[25489] <= r_data[25488];
                
                r_data[25490] <= r_data[25489];
                
                r_data[25491] <= r_data[25490];
                
                r_data[25492] <= r_data[25491];
                
                r_data[25493] <= r_data[25492];
                
                r_data[25494] <= r_data[25493];
                
                r_data[25495] <= r_data[25494];
                
                r_data[25496] <= r_data[25495];
                
                r_data[25497] <= r_data[25496];
                
                r_data[25498] <= r_data[25497];
                
                r_data[25499] <= r_data[25498];
                
                r_data[25500] <= r_data[25499];
                
                r_data[25501] <= r_data[25500];
                
                r_data[25502] <= r_data[25501];
                
                r_data[25503] <= r_data[25502];
                
                r_data[25504] <= r_data[25503];
                
                r_data[25505] <= r_data[25504];
                
                r_data[25506] <= r_data[25505];
                
                r_data[25507] <= r_data[25506];
                
                r_data[25508] <= r_data[25507];
                
                r_data[25509] <= r_data[25508];
                
                r_data[25510] <= r_data[25509];
                
                r_data[25511] <= r_data[25510];
                
                r_data[25512] <= r_data[25511];
                
                r_data[25513] <= r_data[25512];
                
                r_data[25514] <= r_data[25513];
                
                r_data[25515] <= r_data[25514];
                
                r_data[25516] <= r_data[25515];
                
                r_data[25517] <= r_data[25516];
                
                r_data[25518] <= r_data[25517];
                
                r_data[25519] <= r_data[25518];
                
                r_data[25520] <= r_data[25519];
                
                r_data[25521] <= r_data[25520];
                
                r_data[25522] <= r_data[25521];
                
                r_data[25523] <= r_data[25522];
                
                r_data[25524] <= r_data[25523];
                
                r_data[25525] <= r_data[25524];
                
                r_data[25526] <= r_data[25525];
                
                r_data[25527] <= r_data[25526];
                
                r_data[25528] <= r_data[25527];
                
                r_data[25529] <= r_data[25528];
                
                r_data[25530] <= r_data[25529];
                
                r_data[25531] <= r_data[25530];
                
                r_data[25532] <= r_data[25531];
                
                r_data[25533] <= r_data[25532];
                
                r_data[25534] <= r_data[25533];
                
                r_data[25535] <= r_data[25534];
                
                r_data[25536] <= r_data[25535];
                
                r_data[25537] <= r_data[25536];
                
                r_data[25538] <= r_data[25537];
                
                r_data[25539] <= r_data[25538];
                
                r_data[25540] <= r_data[25539];
                
                r_data[25541] <= r_data[25540];
                
                r_data[25542] <= r_data[25541];
                
                r_data[25543] <= r_data[25542];
                
                r_data[25544] <= r_data[25543];
                
                r_data[25545] <= r_data[25544];
                
                r_data[25546] <= r_data[25545];
                
                r_data[25547] <= r_data[25546];
                
                r_data[25548] <= r_data[25547];
                
                r_data[25549] <= r_data[25548];
                
                r_data[25550] <= r_data[25549];
                
                r_data[25551] <= r_data[25550];
                
                r_data[25552] <= r_data[25551];
                
                r_data[25553] <= r_data[25552];
                
                r_data[25554] <= r_data[25553];
                
                r_data[25555] <= r_data[25554];
                
                r_data[25556] <= r_data[25555];
                
                r_data[25557] <= r_data[25556];
                
                r_data[25558] <= r_data[25557];
                
                r_data[25559] <= r_data[25558];
                
                r_data[25560] <= r_data[25559];
                
                r_data[25561] <= r_data[25560];
                
                r_data[25562] <= r_data[25561];
                
                r_data[25563] <= r_data[25562];
                
                r_data[25564] <= r_data[25563];
                
                r_data[25565] <= r_data[25564];
                
                r_data[25566] <= r_data[25565];
                
                r_data[25567] <= r_data[25566];
                
                r_data[25568] <= r_data[25567];
                
                r_data[25569] <= r_data[25568];
                
                r_data[25570] <= r_data[25569];
                
                r_data[25571] <= r_data[25570];
                
                r_data[25572] <= r_data[25571];
                
                r_data[25573] <= r_data[25572];
                
                r_data[25574] <= r_data[25573];
                
                r_data[25575] <= r_data[25574];
                
                r_data[25576] <= r_data[25575];
                
                r_data[25577] <= r_data[25576];
                
                r_data[25578] <= r_data[25577];
                
                r_data[25579] <= r_data[25578];
                
                r_data[25580] <= r_data[25579];
                
                r_data[25581] <= r_data[25580];
                
                r_data[25582] <= r_data[25581];
                
                r_data[25583] <= r_data[25582];
                
                r_data[25584] <= r_data[25583];
                
                r_data[25585] <= r_data[25584];
                
                r_data[25586] <= r_data[25585];
                
                r_data[25587] <= r_data[25586];
                
                r_data[25588] <= r_data[25587];
                
                r_data[25589] <= r_data[25588];
                
                r_data[25590] <= r_data[25589];
                
                r_data[25591] <= r_data[25590];
                
                r_data[25592] <= r_data[25591];
                
                r_data[25593] <= r_data[25592];
                
                r_data[25594] <= r_data[25593];
                
                r_data[25595] <= r_data[25594];
                
                r_data[25596] <= r_data[25595];
                
                r_data[25597] <= r_data[25596];
                
                r_data[25598] <= r_data[25597];
                
                r_data[25599] <= r_data[25598];
                
                r_data[25600] <= r_data[25599];
                
                r_data[25601] <= r_data[25600];
                
                r_data[25602] <= r_data[25601];
                
                r_data[25603] <= r_data[25602];
                
                r_data[25604] <= r_data[25603];
                
                r_data[25605] <= r_data[25604];
                
                r_data[25606] <= r_data[25605];
                
                r_data[25607] <= r_data[25606];
                
                r_data[25608] <= r_data[25607];
                
                r_data[25609] <= r_data[25608];
                
                r_data[25610] <= r_data[25609];
                
                r_data[25611] <= r_data[25610];
                
                r_data[25612] <= r_data[25611];
                
                r_data[25613] <= r_data[25612];
                
                r_data[25614] <= r_data[25613];
                
                r_data[25615] <= r_data[25614];
                
                r_data[25616] <= r_data[25615];
                
                r_data[25617] <= r_data[25616];
                
                r_data[25618] <= r_data[25617];
                
                r_data[25619] <= r_data[25618];
                
                r_data[25620] <= r_data[25619];
                
                r_data[25621] <= r_data[25620];
                
                r_data[25622] <= r_data[25621];
                
                r_data[25623] <= r_data[25622];
                
                r_data[25624] <= r_data[25623];
                
                r_data[25625] <= r_data[25624];
                
                r_data[25626] <= r_data[25625];
                
                r_data[25627] <= r_data[25626];
                
                r_data[25628] <= r_data[25627];
                
                r_data[25629] <= r_data[25628];
                
                r_data[25630] <= r_data[25629];
                
                r_data[25631] <= r_data[25630];
                
                r_data[25632] <= r_data[25631];
                
                r_data[25633] <= r_data[25632];
                
                r_data[25634] <= r_data[25633];
                
                r_data[25635] <= r_data[25634];
                
                r_data[25636] <= r_data[25635];
                
                r_data[25637] <= r_data[25636];
                
                r_data[25638] <= r_data[25637];
                
                r_data[25639] <= r_data[25638];
                
                r_data[25640] <= r_data[25639];
                
                r_data[25641] <= r_data[25640];
                
                r_data[25642] <= r_data[25641];
                
                r_data[25643] <= r_data[25642];
                
                r_data[25644] <= r_data[25643];
                
                r_data[25645] <= r_data[25644];
                
                r_data[25646] <= r_data[25645];
                
                r_data[25647] <= r_data[25646];
                
                r_data[25648] <= r_data[25647];
                
                r_data[25649] <= r_data[25648];
                
                r_data[25650] <= r_data[25649];
                
                r_data[25651] <= r_data[25650];
                
                r_data[25652] <= r_data[25651];
                
                r_data[25653] <= r_data[25652];
                
                r_data[25654] <= r_data[25653];
                
                r_data[25655] <= r_data[25654];
                
                r_data[25656] <= r_data[25655];
                
                r_data[25657] <= r_data[25656];
                
                r_data[25658] <= r_data[25657];
                
                r_data[25659] <= r_data[25658];
                
                r_data[25660] <= r_data[25659];
                
                r_data[25661] <= r_data[25660];
                
                r_data[25662] <= r_data[25661];
                
                r_data[25663] <= r_data[25662];
                
                r_data[25664] <= r_data[25663];
                
                r_data[25665] <= r_data[25664];
                
                r_data[25666] <= r_data[25665];
                
                r_data[25667] <= r_data[25666];
                
                r_data[25668] <= r_data[25667];
                
                r_data[25669] <= r_data[25668];
                
                r_data[25670] <= r_data[25669];
                
                r_data[25671] <= r_data[25670];
                
                r_data[25672] <= r_data[25671];
                
                r_data[25673] <= r_data[25672];
                
                r_data[25674] <= r_data[25673];
                
                r_data[25675] <= r_data[25674];
                
                r_data[25676] <= r_data[25675];
                
                r_data[25677] <= r_data[25676];
                
                r_data[25678] <= r_data[25677];
                
                r_data[25679] <= r_data[25678];
                
                r_data[25680] <= r_data[25679];
                
                r_data[25681] <= r_data[25680];
                
                r_data[25682] <= r_data[25681];
                
                r_data[25683] <= r_data[25682];
                
                r_data[25684] <= r_data[25683];
                
                r_data[25685] <= r_data[25684];
                
                r_data[25686] <= r_data[25685];
                
                r_data[25687] <= r_data[25686];
                
                r_data[25688] <= r_data[25687];
                
                r_data[25689] <= r_data[25688];
                
                r_data[25690] <= r_data[25689];
                
                r_data[25691] <= r_data[25690];
                
                r_data[25692] <= r_data[25691];
                
                r_data[25693] <= r_data[25692];
                
                r_data[25694] <= r_data[25693];
                
                r_data[25695] <= r_data[25694];
                
                r_data[25696] <= r_data[25695];
                
                r_data[25697] <= r_data[25696];
                
                r_data[25698] <= r_data[25697];
                
                r_data[25699] <= r_data[25698];
                
                r_data[25700] <= r_data[25699];
                
                r_data[25701] <= r_data[25700];
                
                r_data[25702] <= r_data[25701];
                
                r_data[25703] <= r_data[25702];
                
                r_data[25704] <= r_data[25703];
                
                r_data[25705] <= r_data[25704];
                
                r_data[25706] <= r_data[25705];
                
                r_data[25707] <= r_data[25706];
                
                r_data[25708] <= r_data[25707];
                
                r_data[25709] <= r_data[25708];
                
                r_data[25710] <= r_data[25709];
                
                r_data[25711] <= r_data[25710];
                
                r_data[25712] <= r_data[25711];
                
                r_data[25713] <= r_data[25712];
                
                r_data[25714] <= r_data[25713];
                
                r_data[25715] <= r_data[25714];
                
                r_data[25716] <= r_data[25715];
                
                r_data[25717] <= r_data[25716];
                
                r_data[25718] <= r_data[25717];
                
                r_data[25719] <= r_data[25718];
                
                r_data[25720] <= r_data[25719];
                
                r_data[25721] <= r_data[25720];
                
                r_data[25722] <= r_data[25721];
                
                r_data[25723] <= r_data[25722];
                
                r_data[25724] <= r_data[25723];
                
                r_data[25725] <= r_data[25724];
                
                r_data[25726] <= r_data[25725];
                
                r_data[25727] <= r_data[25726];
                
                r_data[25728] <= r_data[25727];
                
                r_data[25729] <= r_data[25728];
                
                r_data[25730] <= r_data[25729];
                
                r_data[25731] <= r_data[25730];
                
                r_data[25732] <= r_data[25731];
                
                r_data[25733] <= r_data[25732];
                
                r_data[25734] <= r_data[25733];
                
                r_data[25735] <= r_data[25734];
                
                r_data[25736] <= r_data[25735];
                
                r_data[25737] <= r_data[25736];
                
                r_data[25738] <= r_data[25737];
                
                r_data[25739] <= r_data[25738];
                
                r_data[25740] <= r_data[25739];
                
                r_data[25741] <= r_data[25740];
                
                r_data[25742] <= r_data[25741];
                
                r_data[25743] <= r_data[25742];
                
                r_data[25744] <= r_data[25743];
                
                r_data[25745] <= r_data[25744];
                
                r_data[25746] <= r_data[25745];
                
                r_data[25747] <= r_data[25746];
                
                r_data[25748] <= r_data[25747];
                
                r_data[25749] <= r_data[25748];
                
                r_data[25750] <= r_data[25749];
                
                r_data[25751] <= r_data[25750];
                
                r_data[25752] <= r_data[25751];
                
                r_data[25753] <= r_data[25752];
                
                r_data[25754] <= r_data[25753];
                
                r_data[25755] <= r_data[25754];
                
                r_data[25756] <= r_data[25755];
                
                r_data[25757] <= r_data[25756];
                
                r_data[25758] <= r_data[25757];
                
                r_data[25759] <= r_data[25758];
                
                r_data[25760] <= r_data[25759];
                
                r_data[25761] <= r_data[25760];
                
                r_data[25762] <= r_data[25761];
                
                r_data[25763] <= r_data[25762];
                
                r_data[25764] <= r_data[25763];
                
                r_data[25765] <= r_data[25764];
                
                r_data[25766] <= r_data[25765];
                
                r_data[25767] <= r_data[25766];
                
                r_data[25768] <= r_data[25767];
                
                r_data[25769] <= r_data[25768];
                
                r_data[25770] <= r_data[25769];
                
                r_data[25771] <= r_data[25770];
                
                r_data[25772] <= r_data[25771];
                
                r_data[25773] <= r_data[25772];
                
                r_data[25774] <= r_data[25773];
                
                r_data[25775] <= r_data[25774];
                
                r_data[25776] <= r_data[25775];
                
                r_data[25777] <= r_data[25776];
                
                r_data[25778] <= r_data[25777];
                
                r_data[25779] <= r_data[25778];
                
                r_data[25780] <= r_data[25779];
                
                r_data[25781] <= r_data[25780];
                
                r_data[25782] <= r_data[25781];
                
                r_data[25783] <= r_data[25782];
                
                r_data[25784] <= r_data[25783];
                
                r_data[25785] <= r_data[25784];
                
                r_data[25786] <= r_data[25785];
                
                r_data[25787] <= r_data[25786];
                
                r_data[25788] <= r_data[25787];
                
                r_data[25789] <= r_data[25788];
                
                r_data[25790] <= r_data[25789];
                
                r_data[25791] <= r_data[25790];
                
                r_data[25792] <= r_data[25791];
                
                r_data[25793] <= r_data[25792];
                
                r_data[25794] <= r_data[25793];
                
                r_data[25795] <= r_data[25794];
                
                r_data[25796] <= r_data[25795];
                
                r_data[25797] <= r_data[25796];
                
                r_data[25798] <= r_data[25797];
                
                r_data[25799] <= r_data[25798];
                
                r_data[25800] <= r_data[25799];
                
                r_data[25801] <= r_data[25800];
                
                r_data[25802] <= r_data[25801];
                
                r_data[25803] <= r_data[25802];
                
                r_data[25804] <= r_data[25803];
                
                r_data[25805] <= r_data[25804];
                
                r_data[25806] <= r_data[25805];
                
                r_data[25807] <= r_data[25806];
                
                r_data[25808] <= r_data[25807];
                
                r_data[25809] <= r_data[25808];
                
                r_data[25810] <= r_data[25809];
                
                r_data[25811] <= r_data[25810];
                
                r_data[25812] <= r_data[25811];
                
                r_data[25813] <= r_data[25812];
                
                r_data[25814] <= r_data[25813];
                
                r_data[25815] <= r_data[25814];
                
                r_data[25816] <= r_data[25815];
                
                r_data[25817] <= r_data[25816];
                
                r_data[25818] <= r_data[25817];
                
                r_data[25819] <= r_data[25818];
                
                r_data[25820] <= r_data[25819];
                
                r_data[25821] <= r_data[25820];
                
                r_data[25822] <= r_data[25821];
                
                r_data[25823] <= r_data[25822];
                
                r_data[25824] <= r_data[25823];
                
                r_data[25825] <= r_data[25824];
                
                r_data[25826] <= r_data[25825];
                
                r_data[25827] <= r_data[25826];
                
                r_data[25828] <= r_data[25827];
                
                r_data[25829] <= r_data[25828];
                
                r_data[25830] <= r_data[25829];
                
                r_data[25831] <= r_data[25830];
                
                r_data[25832] <= r_data[25831];
                
                r_data[25833] <= r_data[25832];
                
                r_data[25834] <= r_data[25833];
                
                r_data[25835] <= r_data[25834];
                
                r_data[25836] <= r_data[25835];
                
                r_data[25837] <= r_data[25836];
                
                r_data[25838] <= r_data[25837];
                
                r_data[25839] <= r_data[25838];
                
                r_data[25840] <= r_data[25839];
                
                r_data[25841] <= r_data[25840];
                
                r_data[25842] <= r_data[25841];
                
                r_data[25843] <= r_data[25842];
                
                r_data[25844] <= r_data[25843];
                
                r_data[25845] <= r_data[25844];
                
                r_data[25846] <= r_data[25845];
                
                r_data[25847] <= r_data[25846];
                
                r_data[25848] <= r_data[25847];
                
                r_data[25849] <= r_data[25848];
                
                r_data[25850] <= r_data[25849];
                
                r_data[25851] <= r_data[25850];
                
                r_data[25852] <= r_data[25851];
                
                r_data[25853] <= r_data[25852];
                
                r_data[25854] <= r_data[25853];
                
                r_data[25855] <= r_data[25854];
                
                r_data[25856] <= r_data[25855];
                
                r_data[25857] <= r_data[25856];
                
                r_data[25858] <= r_data[25857];
                
                r_data[25859] <= r_data[25858];
                
                r_data[25860] <= r_data[25859];
                
                r_data[25861] <= r_data[25860];
                
                r_data[25862] <= r_data[25861];
                
                r_data[25863] <= r_data[25862];
                
                r_data[25864] <= r_data[25863];
                
                r_data[25865] <= r_data[25864];
                
                r_data[25866] <= r_data[25865];
                
                r_data[25867] <= r_data[25866];
                
                r_data[25868] <= r_data[25867];
                
                r_data[25869] <= r_data[25868];
                
                r_data[25870] <= r_data[25869];
                
                r_data[25871] <= r_data[25870];
                
                r_data[25872] <= r_data[25871];
                
                r_data[25873] <= r_data[25872];
                
                r_data[25874] <= r_data[25873];
                
                r_data[25875] <= r_data[25874];
                
                r_data[25876] <= r_data[25875];
                
                r_data[25877] <= r_data[25876];
                
                r_data[25878] <= r_data[25877];
                
                r_data[25879] <= r_data[25878];
                
                r_data[25880] <= r_data[25879];
                
                r_data[25881] <= r_data[25880];
                
                r_data[25882] <= r_data[25881];
                
                r_data[25883] <= r_data[25882];
                
                r_data[25884] <= r_data[25883];
                
                r_data[25885] <= r_data[25884];
                
                r_data[25886] <= r_data[25885];
                
                r_data[25887] <= r_data[25886];
                
                r_data[25888] <= r_data[25887];
                
                r_data[25889] <= r_data[25888];
                
                r_data[25890] <= r_data[25889];
                
                r_data[25891] <= r_data[25890];
                
                r_data[25892] <= r_data[25891];
                
                r_data[25893] <= r_data[25892];
                
                r_data[25894] <= r_data[25893];
                
                r_data[25895] <= r_data[25894];
                
                r_data[25896] <= r_data[25895];
                
                r_data[25897] <= r_data[25896];
                
                r_data[25898] <= r_data[25897];
                
                r_data[25899] <= r_data[25898];
                
                r_data[25900] <= r_data[25899];
                
                r_data[25901] <= r_data[25900];
                
                r_data[25902] <= r_data[25901];
                
                r_data[25903] <= r_data[25902];
                
                r_data[25904] <= r_data[25903];
                
                r_data[25905] <= r_data[25904];
                
                r_data[25906] <= r_data[25905];
                
                r_data[25907] <= r_data[25906];
                
                r_data[25908] <= r_data[25907];
                
                r_data[25909] <= r_data[25908];
                
                r_data[25910] <= r_data[25909];
                
                r_data[25911] <= r_data[25910];
                
                r_data[25912] <= r_data[25911];
                
                r_data[25913] <= r_data[25912];
                
                r_data[25914] <= r_data[25913];
                
                r_data[25915] <= r_data[25914];
                
                r_data[25916] <= r_data[25915];
                
                r_data[25917] <= r_data[25916];
                
                r_data[25918] <= r_data[25917];
                
                r_data[25919] <= r_data[25918];
                
                r_data[25920] <= r_data[25919];
                
                r_data[25921] <= r_data[25920];
                
                r_data[25922] <= r_data[25921];
                
                r_data[25923] <= r_data[25922];
                
                r_data[25924] <= r_data[25923];
                
                r_data[25925] <= r_data[25924];
                
                r_data[25926] <= r_data[25925];
                
                r_data[25927] <= r_data[25926];
                
                r_data[25928] <= r_data[25927];
                
                r_data[25929] <= r_data[25928];
                
                r_data[25930] <= r_data[25929];
                
                r_data[25931] <= r_data[25930];
                
                r_data[25932] <= r_data[25931];
                
                r_data[25933] <= r_data[25932];
                
                r_data[25934] <= r_data[25933];
                
                r_data[25935] <= r_data[25934];
                
                r_data[25936] <= r_data[25935];
                
                r_data[25937] <= r_data[25936];
                
                r_data[25938] <= r_data[25937];
                
                r_data[25939] <= r_data[25938];
                
                r_data[25940] <= r_data[25939];
                
                r_data[25941] <= r_data[25940];
                
                r_data[25942] <= r_data[25941];
                
                r_data[25943] <= r_data[25942];
                
                r_data[25944] <= r_data[25943];
                
                r_data[25945] <= r_data[25944];
                
                r_data[25946] <= r_data[25945];
                
                r_data[25947] <= r_data[25946];
                
                r_data[25948] <= r_data[25947];
                
                r_data[25949] <= r_data[25948];
                
                r_data[25950] <= r_data[25949];
                
                r_data[25951] <= r_data[25950];
                
                r_data[25952] <= r_data[25951];
                
                r_data[25953] <= r_data[25952];
                
                r_data[25954] <= r_data[25953];
                
                r_data[25955] <= r_data[25954];
                
                r_data[25956] <= r_data[25955];
                
                r_data[25957] <= r_data[25956];
                
                r_data[25958] <= r_data[25957];
                
                r_data[25959] <= r_data[25958];
                
                r_data[25960] <= r_data[25959];
                
                r_data[25961] <= r_data[25960];
                
                r_data[25962] <= r_data[25961];
                
                r_data[25963] <= r_data[25962];
                
                r_data[25964] <= r_data[25963];
                
                r_data[25965] <= r_data[25964];
                
                r_data[25966] <= r_data[25965];
                
                r_data[25967] <= r_data[25966];
                
                r_data[25968] <= r_data[25967];
                
                r_data[25969] <= r_data[25968];
                
                r_data[25970] <= r_data[25969];
                
                r_data[25971] <= r_data[25970];
                
                r_data[25972] <= r_data[25971];
                
                r_data[25973] <= r_data[25972];
                
                r_data[25974] <= r_data[25973];
                
                r_data[25975] <= r_data[25974];
                
                r_data[25976] <= r_data[25975];
                
                r_data[25977] <= r_data[25976];
                
                r_data[25978] <= r_data[25977];
                
                r_data[25979] <= r_data[25978];
                
                r_data[25980] <= r_data[25979];
                
                r_data[25981] <= r_data[25980];
                
                r_data[25982] <= r_data[25981];
                
                r_data[25983] <= r_data[25982];
                
                r_data[25984] <= r_data[25983];
                
                r_data[25985] <= r_data[25984];
                
                r_data[25986] <= r_data[25985];
                
                r_data[25987] <= r_data[25986];
                
                r_data[25988] <= r_data[25987];
                
                r_data[25989] <= r_data[25988];
                
                r_data[25990] <= r_data[25989];
                
                r_data[25991] <= r_data[25990];
                
                r_data[25992] <= r_data[25991];
                
                r_data[25993] <= r_data[25992];
                
                r_data[25994] <= r_data[25993];
                
                r_data[25995] <= r_data[25994];
                
                r_data[25996] <= r_data[25995];
                
                r_data[25997] <= r_data[25996];
                
                r_data[25998] <= r_data[25997];
                
                r_data[25999] <= r_data[25998];
                
                r_data[26000] <= r_data[25999];
                
                r_data[26001] <= r_data[26000];
                
                r_data[26002] <= r_data[26001];
                
                r_data[26003] <= r_data[26002];
                
                r_data[26004] <= r_data[26003];
                
                r_data[26005] <= r_data[26004];
                
                r_data[26006] <= r_data[26005];
                
                r_data[26007] <= r_data[26006];
                
                r_data[26008] <= r_data[26007];
                
                r_data[26009] <= r_data[26008];
                
                r_data[26010] <= r_data[26009];
                
                r_data[26011] <= r_data[26010];
                
                r_data[26012] <= r_data[26011];
                
                r_data[26013] <= r_data[26012];
                
                r_data[26014] <= r_data[26013];
                
                r_data[26015] <= r_data[26014];
                
                r_data[26016] <= r_data[26015];
                
                r_data[26017] <= r_data[26016];
                
                r_data[26018] <= r_data[26017];
                
                r_data[26019] <= r_data[26018];
                
                r_data[26020] <= r_data[26019];
                
                r_data[26021] <= r_data[26020];
                
                r_data[26022] <= r_data[26021];
                
                r_data[26023] <= r_data[26022];
                
                r_data[26024] <= r_data[26023];
                
                r_data[26025] <= r_data[26024];
                
                r_data[26026] <= r_data[26025];
                
                r_data[26027] <= r_data[26026];
                
                r_data[26028] <= r_data[26027];
                
                r_data[26029] <= r_data[26028];
                
                r_data[26030] <= r_data[26029];
                
                r_data[26031] <= r_data[26030];
                
                r_data[26032] <= r_data[26031];
                
                r_data[26033] <= r_data[26032];
                
                r_data[26034] <= r_data[26033];
                
                r_data[26035] <= r_data[26034];
                
                r_data[26036] <= r_data[26035];
                
                r_data[26037] <= r_data[26036];
                
                r_data[26038] <= r_data[26037];
                
                r_data[26039] <= r_data[26038];
                
                r_data[26040] <= r_data[26039];
                
                r_data[26041] <= r_data[26040];
                
                r_data[26042] <= r_data[26041];
                
                r_data[26043] <= r_data[26042];
                
                r_data[26044] <= r_data[26043];
                
                r_data[26045] <= r_data[26044];
                
                r_data[26046] <= r_data[26045];
                
                r_data[26047] <= r_data[26046];
                
                r_data[26048] <= r_data[26047];
                
                r_data[26049] <= r_data[26048];
                
                r_data[26050] <= r_data[26049];
                
                r_data[26051] <= r_data[26050];
                
                r_data[26052] <= r_data[26051];
                
                r_data[26053] <= r_data[26052];
                
                r_data[26054] <= r_data[26053];
                
                r_data[26055] <= r_data[26054];
                
                r_data[26056] <= r_data[26055];
                
                r_data[26057] <= r_data[26056];
                
                r_data[26058] <= r_data[26057];
                
                r_data[26059] <= r_data[26058];
                
                r_data[26060] <= r_data[26059];
                
                r_data[26061] <= r_data[26060];
                
                r_data[26062] <= r_data[26061];
                
                r_data[26063] <= r_data[26062];
                
                r_data[26064] <= r_data[26063];
                
                r_data[26065] <= r_data[26064];
                
                r_data[26066] <= r_data[26065];
                
                r_data[26067] <= r_data[26066];
                
                r_data[26068] <= r_data[26067];
                
                r_data[26069] <= r_data[26068];
                
                r_data[26070] <= r_data[26069];
                
                r_data[26071] <= r_data[26070];
                
                r_data[26072] <= r_data[26071];
                
                r_data[26073] <= r_data[26072];
                
                r_data[26074] <= r_data[26073];
                
                r_data[26075] <= r_data[26074];
                
                r_data[26076] <= r_data[26075];
                
                r_data[26077] <= r_data[26076];
                
                r_data[26078] <= r_data[26077];
                
                r_data[26079] <= r_data[26078];
                
                r_data[26080] <= r_data[26079];
                
                r_data[26081] <= r_data[26080];
                
                r_data[26082] <= r_data[26081];
                
                r_data[26083] <= r_data[26082];
                
                r_data[26084] <= r_data[26083];
                
                r_data[26085] <= r_data[26084];
                
                r_data[26086] <= r_data[26085];
                
                r_data[26087] <= r_data[26086];
                
                r_data[26088] <= r_data[26087];
                
                r_data[26089] <= r_data[26088];
                
                r_data[26090] <= r_data[26089];
                
                r_data[26091] <= r_data[26090];
                
                r_data[26092] <= r_data[26091];
                
                r_data[26093] <= r_data[26092];
                
                r_data[26094] <= r_data[26093];
                
                r_data[26095] <= r_data[26094];
                
                r_data[26096] <= r_data[26095];
                
                r_data[26097] <= r_data[26096];
                
                r_data[26098] <= r_data[26097];
                
                r_data[26099] <= r_data[26098];
                
                r_data[26100] <= r_data[26099];
                
                r_data[26101] <= r_data[26100];
                
                r_data[26102] <= r_data[26101];
                
                r_data[26103] <= r_data[26102];
                
                r_data[26104] <= r_data[26103];
                
                r_data[26105] <= r_data[26104];
                
                r_data[26106] <= r_data[26105];
                
                r_data[26107] <= r_data[26106];
                
                r_data[26108] <= r_data[26107];
                
                r_data[26109] <= r_data[26108];
                
                r_data[26110] <= r_data[26109];
                
                r_data[26111] <= r_data[26110];
                
                r_data[26112] <= r_data[26111];
                
                r_data[26113] <= r_data[26112];
                
                r_data[26114] <= r_data[26113];
                
                r_data[26115] <= r_data[26114];
                
                r_data[26116] <= r_data[26115];
                
                r_data[26117] <= r_data[26116];
                
                r_data[26118] <= r_data[26117];
                
                r_data[26119] <= r_data[26118];
                
                r_data[26120] <= r_data[26119];
                
                r_data[26121] <= r_data[26120];
                
                r_data[26122] <= r_data[26121];
                
                r_data[26123] <= r_data[26122];
                
                r_data[26124] <= r_data[26123];
                
                r_data[26125] <= r_data[26124];
                
                r_data[26126] <= r_data[26125];
                
                r_data[26127] <= r_data[26126];
                
                r_data[26128] <= r_data[26127];
                
                r_data[26129] <= r_data[26128];
                
                r_data[26130] <= r_data[26129];
                
                r_data[26131] <= r_data[26130];
                
                r_data[26132] <= r_data[26131];
                
                r_data[26133] <= r_data[26132];
                
                r_data[26134] <= r_data[26133];
                
                r_data[26135] <= r_data[26134];
                
                r_data[26136] <= r_data[26135];
                
                r_data[26137] <= r_data[26136];
                
                r_data[26138] <= r_data[26137];
                
                r_data[26139] <= r_data[26138];
                
                r_data[26140] <= r_data[26139];
                
                r_data[26141] <= r_data[26140];
                
                r_data[26142] <= r_data[26141];
                
                r_data[26143] <= r_data[26142];
                
                r_data[26144] <= r_data[26143];
                
                r_data[26145] <= r_data[26144];
                
                r_data[26146] <= r_data[26145];
                
                r_data[26147] <= r_data[26146];
                
                r_data[26148] <= r_data[26147];
                
                r_data[26149] <= r_data[26148];
                
                r_data[26150] <= r_data[26149];
                
                r_data[26151] <= r_data[26150];
                
                r_data[26152] <= r_data[26151];
                
                r_data[26153] <= r_data[26152];
                
                r_data[26154] <= r_data[26153];
                
                r_data[26155] <= r_data[26154];
                
                r_data[26156] <= r_data[26155];
                
                r_data[26157] <= r_data[26156];
                
                r_data[26158] <= r_data[26157];
                
                r_data[26159] <= r_data[26158];
                
                r_data[26160] <= r_data[26159];
                
                r_data[26161] <= r_data[26160];
                
                r_data[26162] <= r_data[26161];
                
                r_data[26163] <= r_data[26162];
                
                r_data[26164] <= r_data[26163];
                
                r_data[26165] <= r_data[26164];
                
                r_data[26166] <= r_data[26165];
                
                r_data[26167] <= r_data[26166];
                
                r_data[26168] <= r_data[26167];
                
                r_data[26169] <= r_data[26168];
                
                r_data[26170] <= r_data[26169];
                
                r_data[26171] <= r_data[26170];
                
                r_data[26172] <= r_data[26171];
                
                r_data[26173] <= r_data[26172];
                
                r_data[26174] <= r_data[26173];
                
                r_data[26175] <= r_data[26174];
                
                r_data[26176] <= r_data[26175];
                
                r_data[26177] <= r_data[26176];
                
                r_data[26178] <= r_data[26177];
                
                r_data[26179] <= r_data[26178];
                
                r_data[26180] <= r_data[26179];
                
                r_data[26181] <= r_data[26180];
                
                r_data[26182] <= r_data[26181];
                
                r_data[26183] <= r_data[26182];
                
                r_data[26184] <= r_data[26183];
                
                r_data[26185] <= r_data[26184];
                
                r_data[26186] <= r_data[26185];
                
                r_data[26187] <= r_data[26186];
                
                r_data[26188] <= r_data[26187];
                
                r_data[26189] <= r_data[26188];
                
                r_data[26190] <= r_data[26189];
                
                r_data[26191] <= r_data[26190];
                
                r_data[26192] <= r_data[26191];
                
                r_data[26193] <= r_data[26192];
                
                r_data[26194] <= r_data[26193];
                
                r_data[26195] <= r_data[26194];
                
                r_data[26196] <= r_data[26195];
                
                r_data[26197] <= r_data[26196];
                
                r_data[26198] <= r_data[26197];
                
                r_data[26199] <= r_data[26198];
                
                r_data[26200] <= r_data[26199];
                
                r_data[26201] <= r_data[26200];
                
                r_data[26202] <= r_data[26201];
                
                r_data[26203] <= r_data[26202];
                
                r_data[26204] <= r_data[26203];
                
                r_data[26205] <= r_data[26204];
                
                r_data[26206] <= r_data[26205];
                
                r_data[26207] <= r_data[26206];
                
                r_data[26208] <= r_data[26207];
                
                r_data[26209] <= r_data[26208];
                
                r_data[26210] <= r_data[26209];
                
                r_data[26211] <= r_data[26210];
                
                r_data[26212] <= r_data[26211];
                
                r_data[26213] <= r_data[26212];
                
                r_data[26214] <= r_data[26213];
                
                r_data[26215] <= r_data[26214];
                
                r_data[26216] <= r_data[26215];
                
                r_data[26217] <= r_data[26216];
                
                r_data[26218] <= r_data[26217];
                
                r_data[26219] <= r_data[26218];
                
                r_data[26220] <= r_data[26219];
                
                r_data[26221] <= r_data[26220];
                
                r_data[26222] <= r_data[26221];
                
                r_data[26223] <= r_data[26222];
                
                r_data[26224] <= r_data[26223];
                
                r_data[26225] <= r_data[26224];
                
                r_data[26226] <= r_data[26225];
                
                r_data[26227] <= r_data[26226];
                
                r_data[26228] <= r_data[26227];
                
                r_data[26229] <= r_data[26228];
                
                r_data[26230] <= r_data[26229];
                
                r_data[26231] <= r_data[26230];
                
                r_data[26232] <= r_data[26231];
                
                r_data[26233] <= r_data[26232];
                
                r_data[26234] <= r_data[26233];
                
                r_data[26235] <= r_data[26234];
                
                r_data[26236] <= r_data[26235];
                
                r_data[26237] <= r_data[26236];
                
                r_data[26238] <= r_data[26237];
                
                r_data[26239] <= r_data[26238];
                
                r_data[26240] <= r_data[26239];
                
                r_data[26241] <= r_data[26240];
                
                r_data[26242] <= r_data[26241];
                
                r_data[26243] <= r_data[26242];
                
                r_data[26244] <= r_data[26243];
                
                r_data[26245] <= r_data[26244];
                
                r_data[26246] <= r_data[26245];
                
                r_data[26247] <= r_data[26246];
                
                r_data[26248] <= r_data[26247];
                
                r_data[26249] <= r_data[26248];
                
                r_data[26250] <= r_data[26249];
                
                r_data[26251] <= r_data[26250];
                
                r_data[26252] <= r_data[26251];
                
                r_data[26253] <= r_data[26252];
                
                r_data[26254] <= r_data[26253];
                
                r_data[26255] <= r_data[26254];
                
                r_data[26256] <= r_data[26255];
                
                r_data[26257] <= r_data[26256];
                
                r_data[26258] <= r_data[26257];
                
                r_data[26259] <= r_data[26258];
                
                r_data[26260] <= r_data[26259];
                
                r_data[26261] <= r_data[26260];
                
                r_data[26262] <= r_data[26261];
                
                r_data[26263] <= r_data[26262];
                
                r_data[26264] <= r_data[26263];
                
                r_data[26265] <= r_data[26264];
                
                r_data[26266] <= r_data[26265];
                
                r_data[26267] <= r_data[26266];
                
                r_data[26268] <= r_data[26267];
                
                r_data[26269] <= r_data[26268];
                
                r_data[26270] <= r_data[26269];
                
                r_data[26271] <= r_data[26270];
                
                r_data[26272] <= r_data[26271];
                
                r_data[26273] <= r_data[26272];
                
                r_data[26274] <= r_data[26273];
                
                r_data[26275] <= r_data[26274];
                
                r_data[26276] <= r_data[26275];
                
                r_data[26277] <= r_data[26276];
                
                r_data[26278] <= r_data[26277];
                
                r_data[26279] <= r_data[26278];
                
                r_data[26280] <= r_data[26279];
                
                r_data[26281] <= r_data[26280];
                
                r_data[26282] <= r_data[26281];
                
                r_data[26283] <= r_data[26282];
                
                r_data[26284] <= r_data[26283];
                
                r_data[26285] <= r_data[26284];
                
                r_data[26286] <= r_data[26285];
                
                r_data[26287] <= r_data[26286];
                
                r_data[26288] <= r_data[26287];
                
                r_data[26289] <= r_data[26288];
                
                r_data[26290] <= r_data[26289];
                
                r_data[26291] <= r_data[26290];
                
                r_data[26292] <= r_data[26291];
                
                r_data[26293] <= r_data[26292];
                
                r_data[26294] <= r_data[26293];
                
                r_data[26295] <= r_data[26294];
                
                r_data[26296] <= r_data[26295];
                
                r_data[26297] <= r_data[26296];
                
                r_data[26298] <= r_data[26297];
                
                r_data[26299] <= r_data[26298];
                
                r_data[26300] <= r_data[26299];
                
                r_data[26301] <= r_data[26300];
                
                r_data[26302] <= r_data[26301];
                
                r_data[26303] <= r_data[26302];
                
                r_data[26304] <= r_data[26303];
                
                r_data[26305] <= r_data[26304];
                
                r_data[26306] <= r_data[26305];
                
                r_data[26307] <= r_data[26306];
                
                r_data[26308] <= r_data[26307];
                
                r_data[26309] <= r_data[26308];
                
                r_data[26310] <= r_data[26309];
                
                r_data[26311] <= r_data[26310];
                
                r_data[26312] <= r_data[26311];
                
                r_data[26313] <= r_data[26312];
                
                r_data[26314] <= r_data[26313];
                
                r_data[26315] <= r_data[26314];
                
                r_data[26316] <= r_data[26315];
                
                r_data[26317] <= r_data[26316];
                
                r_data[26318] <= r_data[26317];
                
                r_data[26319] <= r_data[26318];
                
                r_data[26320] <= r_data[26319];
                
                r_data[26321] <= r_data[26320];
                
                r_data[26322] <= r_data[26321];
                
                r_data[26323] <= r_data[26322];
                
                r_data[26324] <= r_data[26323];
                
                r_data[26325] <= r_data[26324];
                
                r_data[26326] <= r_data[26325];
                
                r_data[26327] <= r_data[26326];
                
                r_data[26328] <= r_data[26327];
                
                r_data[26329] <= r_data[26328];
                
                r_data[26330] <= r_data[26329];
                
                r_data[26331] <= r_data[26330];
                
                r_data[26332] <= r_data[26331];
                
                r_data[26333] <= r_data[26332];
                
                r_data[26334] <= r_data[26333];
                
                r_data[26335] <= r_data[26334];
                
                r_data[26336] <= r_data[26335];
                
                r_data[26337] <= r_data[26336];
                
                r_data[26338] <= r_data[26337];
                
                r_data[26339] <= r_data[26338];
                
                r_data[26340] <= r_data[26339];
                
                r_data[26341] <= r_data[26340];
                
                r_data[26342] <= r_data[26341];
                
                r_data[26343] <= r_data[26342];
                
                r_data[26344] <= r_data[26343];
                
                r_data[26345] <= r_data[26344];
                
                r_data[26346] <= r_data[26345];
                
                r_data[26347] <= r_data[26346];
                
                r_data[26348] <= r_data[26347];
                
                r_data[26349] <= r_data[26348];
                
                r_data[26350] <= r_data[26349];
                
                r_data[26351] <= r_data[26350];
                
                r_data[26352] <= r_data[26351];
                
                r_data[26353] <= r_data[26352];
                
                r_data[26354] <= r_data[26353];
                
                r_data[26355] <= r_data[26354];
                
                r_data[26356] <= r_data[26355];
                
                r_data[26357] <= r_data[26356];
                
                r_data[26358] <= r_data[26357];
                
                r_data[26359] <= r_data[26358];
                
                r_data[26360] <= r_data[26359];
                
                r_data[26361] <= r_data[26360];
                
                r_data[26362] <= r_data[26361];
                
                r_data[26363] <= r_data[26362];
                
                r_data[26364] <= r_data[26363];
                
                r_data[26365] <= r_data[26364];
                
                r_data[26366] <= r_data[26365];
                
                r_data[26367] <= r_data[26366];
                
                r_data[26368] <= r_data[26367];
                
                r_data[26369] <= r_data[26368];
                
                r_data[26370] <= r_data[26369];
                
                r_data[26371] <= r_data[26370];
                
                r_data[26372] <= r_data[26371];
                
                r_data[26373] <= r_data[26372];
                
                r_data[26374] <= r_data[26373];
                
                r_data[26375] <= r_data[26374];
                
                r_data[26376] <= r_data[26375];
                
                r_data[26377] <= r_data[26376];
                
                r_data[26378] <= r_data[26377];
                
                r_data[26379] <= r_data[26378];
                
                r_data[26380] <= r_data[26379];
                
                r_data[26381] <= r_data[26380];
                
                r_data[26382] <= r_data[26381];
                
                r_data[26383] <= r_data[26382];
                
                r_data[26384] <= r_data[26383];
                
                r_data[26385] <= r_data[26384];
                
                r_data[26386] <= r_data[26385];
                
                r_data[26387] <= r_data[26386];
                
                r_data[26388] <= r_data[26387];
                
                r_data[26389] <= r_data[26388];
                
                r_data[26390] <= r_data[26389];
                
                r_data[26391] <= r_data[26390];
                
                r_data[26392] <= r_data[26391];
                
                r_data[26393] <= r_data[26392];
                
                r_data[26394] <= r_data[26393];
                
                r_data[26395] <= r_data[26394];
                
                r_data[26396] <= r_data[26395];
                
                r_data[26397] <= r_data[26396];
                
                r_data[26398] <= r_data[26397];
                
                r_data[26399] <= r_data[26398];
                
                r_data[26400] <= r_data[26399];
                
                r_data[26401] <= r_data[26400];
                
                r_data[26402] <= r_data[26401];
                
                r_data[26403] <= r_data[26402];
                
                r_data[26404] <= r_data[26403];
                
                r_data[26405] <= r_data[26404];
                
                r_data[26406] <= r_data[26405];
                
                r_data[26407] <= r_data[26406];
                
                r_data[26408] <= r_data[26407];
                
                r_data[26409] <= r_data[26408];
                
                r_data[26410] <= r_data[26409];
                
                r_data[26411] <= r_data[26410];
                
                r_data[26412] <= r_data[26411];
                
                r_data[26413] <= r_data[26412];
                
                r_data[26414] <= r_data[26413];
                
                r_data[26415] <= r_data[26414];
                
                r_data[26416] <= r_data[26415];
                
                r_data[26417] <= r_data[26416];
                
                r_data[26418] <= r_data[26417];
                
                r_data[26419] <= r_data[26418];
                
                r_data[26420] <= r_data[26419];
                
                r_data[26421] <= r_data[26420];
                
                r_data[26422] <= r_data[26421];
                
                r_data[26423] <= r_data[26422];
                
                r_data[26424] <= r_data[26423];
                
                r_data[26425] <= r_data[26424];
                
                r_data[26426] <= r_data[26425];
                
                r_data[26427] <= r_data[26426];
                
                r_data[26428] <= r_data[26427];
                
                r_data[26429] <= r_data[26428];
                
                r_data[26430] <= r_data[26429];
                
                r_data[26431] <= r_data[26430];
                
                r_data[26432] <= r_data[26431];
                
                r_data[26433] <= r_data[26432];
                
                r_data[26434] <= r_data[26433];
                
                r_data[26435] <= r_data[26434];
                
                r_data[26436] <= r_data[26435];
                
                r_data[26437] <= r_data[26436];
                
                r_data[26438] <= r_data[26437];
                
                r_data[26439] <= r_data[26438];
                
                r_data[26440] <= r_data[26439];
                
                r_data[26441] <= r_data[26440];
                
                r_data[26442] <= r_data[26441];
                
                r_data[26443] <= r_data[26442];
                
                r_data[26444] <= r_data[26443];
                
                r_data[26445] <= r_data[26444];
                
                r_data[26446] <= r_data[26445];
                
                r_data[26447] <= r_data[26446];
                
                r_data[26448] <= r_data[26447];
                
                r_data[26449] <= r_data[26448];
                
                r_data[26450] <= r_data[26449];
                
                r_data[26451] <= r_data[26450];
                
                r_data[26452] <= r_data[26451];
                
                r_data[26453] <= r_data[26452];
                
                r_data[26454] <= r_data[26453];
                
                r_data[26455] <= r_data[26454];
                
                r_data[26456] <= r_data[26455];
                
                r_data[26457] <= r_data[26456];
                
                r_data[26458] <= r_data[26457];
                
                r_data[26459] <= r_data[26458];
                
                r_data[26460] <= r_data[26459];
                
                r_data[26461] <= r_data[26460];
                
                r_data[26462] <= r_data[26461];
                
                r_data[26463] <= r_data[26462];
                
                r_data[26464] <= r_data[26463];
                
                r_data[26465] <= r_data[26464];
                
                r_data[26466] <= r_data[26465];
                
                r_data[26467] <= r_data[26466];
                
                r_data[26468] <= r_data[26467];
                
                r_data[26469] <= r_data[26468];
                
                r_data[26470] <= r_data[26469];
                
                r_data[26471] <= r_data[26470];
                
                r_data[26472] <= r_data[26471];
                
                r_data[26473] <= r_data[26472];
                
                r_data[26474] <= r_data[26473];
                
                r_data[26475] <= r_data[26474];
                
                r_data[26476] <= r_data[26475];
                
                r_data[26477] <= r_data[26476];
                
                r_data[26478] <= r_data[26477];
                
                r_data[26479] <= r_data[26478];
                
                r_data[26480] <= r_data[26479];
                
                r_data[26481] <= r_data[26480];
                
                r_data[26482] <= r_data[26481];
                
                r_data[26483] <= r_data[26482];
                
                r_data[26484] <= r_data[26483];
                
                r_data[26485] <= r_data[26484];
                
                r_data[26486] <= r_data[26485];
                
                r_data[26487] <= r_data[26486];
                
                r_data[26488] <= r_data[26487];
                
                r_data[26489] <= r_data[26488];
                
                r_data[26490] <= r_data[26489];
                
                r_data[26491] <= r_data[26490];
                
                r_data[26492] <= r_data[26491];
                
                r_data[26493] <= r_data[26492];
                
                r_data[26494] <= r_data[26493];
                
                r_data[26495] <= r_data[26494];
                
                r_data[26496] <= r_data[26495];
                
                r_data[26497] <= r_data[26496];
                
                r_data[26498] <= r_data[26497];
                
                r_data[26499] <= r_data[26498];
                
                r_data[26500] <= r_data[26499];
                
                r_data[26501] <= r_data[26500];
                
                r_data[26502] <= r_data[26501];
                
                r_data[26503] <= r_data[26502];
                
                r_data[26504] <= r_data[26503];
                
                r_data[26505] <= r_data[26504];
                
                r_data[26506] <= r_data[26505];
                
                r_data[26507] <= r_data[26506];
                
                r_data[26508] <= r_data[26507];
                
                r_data[26509] <= r_data[26508];
                
                r_data[26510] <= r_data[26509];
                
                r_data[26511] <= r_data[26510];
                
                r_data[26512] <= r_data[26511];
                
                r_data[26513] <= r_data[26512];
                
                r_data[26514] <= r_data[26513];
                
                r_data[26515] <= r_data[26514];
                
                r_data[26516] <= r_data[26515];
                
                r_data[26517] <= r_data[26516];
                
                r_data[26518] <= r_data[26517];
                
                r_data[26519] <= r_data[26518];
                
                r_data[26520] <= r_data[26519];
                
                r_data[26521] <= r_data[26520];
                
                r_data[26522] <= r_data[26521];
                
                r_data[26523] <= r_data[26522];
                
                r_data[26524] <= r_data[26523];
                
                r_data[26525] <= r_data[26524];
                
                r_data[26526] <= r_data[26525];
                
                r_data[26527] <= r_data[26526];
                
                r_data[26528] <= r_data[26527];
                
                r_data[26529] <= r_data[26528];
                
                r_data[26530] <= r_data[26529];
                
                r_data[26531] <= r_data[26530];
                
                r_data[26532] <= r_data[26531];
                
                r_data[26533] <= r_data[26532];
                
                r_data[26534] <= r_data[26533];
                
                r_data[26535] <= r_data[26534];
                
                r_data[26536] <= r_data[26535];
                
                r_data[26537] <= r_data[26536];
                
                r_data[26538] <= r_data[26537];
                
                r_data[26539] <= r_data[26538];
                
                r_data[26540] <= r_data[26539];
                
                r_data[26541] <= r_data[26540];
                
                r_data[26542] <= r_data[26541];
                
                r_data[26543] <= r_data[26542];
                
                r_data[26544] <= r_data[26543];
                
                r_data[26545] <= r_data[26544];
                
                r_data[26546] <= r_data[26545];
                
                r_data[26547] <= r_data[26546];
                
                r_data[26548] <= r_data[26547];
                
                r_data[26549] <= r_data[26548];
                
                r_data[26550] <= r_data[26549];
                
                r_data[26551] <= r_data[26550];
                
                r_data[26552] <= r_data[26551];
                
                r_data[26553] <= r_data[26552];
                
                r_data[26554] <= r_data[26553];
                
                r_data[26555] <= r_data[26554];
                
                r_data[26556] <= r_data[26555];
                
                r_data[26557] <= r_data[26556];
                
                r_data[26558] <= r_data[26557];
                
                r_data[26559] <= r_data[26558];
                
                r_data[26560] <= r_data[26559];
                
                r_data[26561] <= r_data[26560];
                
                r_data[26562] <= r_data[26561];
                
                r_data[26563] <= r_data[26562];
                
                r_data[26564] <= r_data[26563];
                
                r_data[26565] <= r_data[26564];
                
                r_data[26566] <= r_data[26565];
                
                r_data[26567] <= r_data[26566];
                
                r_data[26568] <= r_data[26567];
                
                r_data[26569] <= r_data[26568];
                
                r_data[26570] <= r_data[26569];
                
                r_data[26571] <= r_data[26570];
                
                r_data[26572] <= r_data[26571];
                
                r_data[26573] <= r_data[26572];
                
                r_data[26574] <= r_data[26573];
                
                r_data[26575] <= r_data[26574];
                
                r_data[26576] <= r_data[26575];
                
                r_data[26577] <= r_data[26576];
                
                r_data[26578] <= r_data[26577];
                
                r_data[26579] <= r_data[26578];
                
                r_data[26580] <= r_data[26579];
                
                r_data[26581] <= r_data[26580];
                
                r_data[26582] <= r_data[26581];
                
                r_data[26583] <= r_data[26582];
                
                r_data[26584] <= r_data[26583];
                
                r_data[26585] <= r_data[26584];
                
                r_data[26586] <= r_data[26585];
                
                r_data[26587] <= r_data[26586];
                
                r_data[26588] <= r_data[26587];
                
                r_data[26589] <= r_data[26588];
                
                r_data[26590] <= r_data[26589];
                
                r_data[26591] <= r_data[26590];
                
                r_data[26592] <= r_data[26591];
                
                r_data[26593] <= r_data[26592];
                
                r_data[26594] <= r_data[26593];
                
                r_data[26595] <= r_data[26594];
                
                r_data[26596] <= r_data[26595];
                
                r_data[26597] <= r_data[26596];
                
                r_data[26598] <= r_data[26597];
                
                r_data[26599] <= r_data[26598];
                
                r_data[26600] <= r_data[26599];
                
                r_data[26601] <= r_data[26600];
                
                r_data[26602] <= r_data[26601];
                
                r_data[26603] <= r_data[26602];
                
                r_data[26604] <= r_data[26603];
                
                r_data[26605] <= r_data[26604];
                
                r_data[26606] <= r_data[26605];
                
                r_data[26607] <= r_data[26606];
                
                r_data[26608] <= r_data[26607];
                
                r_data[26609] <= r_data[26608];
                
                r_data[26610] <= r_data[26609];
                
                r_data[26611] <= r_data[26610];
                
                r_data[26612] <= r_data[26611];
                
                r_data[26613] <= r_data[26612];
                
                r_data[26614] <= r_data[26613];
                
                r_data[26615] <= r_data[26614];
                
                r_data[26616] <= r_data[26615];
                
                r_data[26617] <= r_data[26616];
                
                r_data[26618] <= r_data[26617];
                
                r_data[26619] <= r_data[26618];
                
                r_data[26620] <= r_data[26619];
                
                r_data[26621] <= r_data[26620];
                
                r_data[26622] <= r_data[26621];
                
                r_data[26623] <= r_data[26622];
                
                r_data[26624] <= r_data[26623];
                
                r_data[26625] <= r_data[26624];
                
                r_data[26626] <= r_data[26625];
                
                r_data[26627] <= r_data[26626];
                
                r_data[26628] <= r_data[26627];
                
                r_data[26629] <= r_data[26628];
                
                r_data[26630] <= r_data[26629];
                
                r_data[26631] <= r_data[26630];
                
                r_data[26632] <= r_data[26631];
                
                r_data[26633] <= r_data[26632];
                
                r_data[26634] <= r_data[26633];
                
                r_data[26635] <= r_data[26634];
                
                r_data[26636] <= r_data[26635];
                
                r_data[26637] <= r_data[26636];
                
                r_data[26638] <= r_data[26637];
                
                r_data[26639] <= r_data[26638];
                
                r_data[26640] <= r_data[26639];
                
                r_data[26641] <= r_data[26640];
                
                r_data[26642] <= r_data[26641];
                
                r_data[26643] <= r_data[26642];
                
                r_data[26644] <= r_data[26643];
                
                r_data[26645] <= r_data[26644];
                
                r_data[26646] <= r_data[26645];
                
                r_data[26647] <= r_data[26646];
                
                r_data[26648] <= r_data[26647];
                
                r_data[26649] <= r_data[26648];
                
                r_data[26650] <= r_data[26649];
                
                r_data[26651] <= r_data[26650];
                
                r_data[26652] <= r_data[26651];
                
                r_data[26653] <= r_data[26652];
                
                r_data[26654] <= r_data[26653];
                
                r_data[26655] <= r_data[26654];
                
                r_data[26656] <= r_data[26655];
                
                r_data[26657] <= r_data[26656];
                
                r_data[26658] <= r_data[26657];
                
                r_data[26659] <= r_data[26658];
                
                r_data[26660] <= r_data[26659];
                
                r_data[26661] <= r_data[26660];
                
                r_data[26662] <= r_data[26661];
                
                r_data[26663] <= r_data[26662];
                
                r_data[26664] <= r_data[26663];
                
                r_data[26665] <= r_data[26664];
                
                r_data[26666] <= r_data[26665];
                
                r_data[26667] <= r_data[26666];
                
                r_data[26668] <= r_data[26667];
                
                r_data[26669] <= r_data[26668];
                
                r_data[26670] <= r_data[26669];
                
                r_data[26671] <= r_data[26670];
                
                r_data[26672] <= r_data[26671];
                
                r_data[26673] <= r_data[26672];
                
                r_data[26674] <= r_data[26673];
                
                r_data[26675] <= r_data[26674];
                
                r_data[26676] <= r_data[26675];
                
                r_data[26677] <= r_data[26676];
                
                r_data[26678] <= r_data[26677];
                
                r_data[26679] <= r_data[26678];
                
                r_data[26680] <= r_data[26679];
                
                r_data[26681] <= r_data[26680];
                
                r_data[26682] <= r_data[26681];
                
                r_data[26683] <= r_data[26682];
                
                r_data[26684] <= r_data[26683];
                
                r_data[26685] <= r_data[26684];
                
                r_data[26686] <= r_data[26685];
                
                r_data[26687] <= r_data[26686];
                
                r_data[26688] <= r_data[26687];
                
                r_data[26689] <= r_data[26688];
                
                r_data[26690] <= r_data[26689];
                
                r_data[26691] <= r_data[26690];
                
                r_data[26692] <= r_data[26691];
                
                r_data[26693] <= r_data[26692];
                
                r_data[26694] <= r_data[26693];
                
                r_data[26695] <= r_data[26694];
                
                r_data[26696] <= r_data[26695];
                
                r_data[26697] <= r_data[26696];
                
                r_data[26698] <= r_data[26697];
                
                r_data[26699] <= r_data[26698];
                
                r_data[26700] <= r_data[26699];
                
                r_data[26701] <= r_data[26700];
                
                r_data[26702] <= r_data[26701];
                
                r_data[26703] <= r_data[26702];
                
                r_data[26704] <= r_data[26703];
                
                r_data[26705] <= r_data[26704];
                
                r_data[26706] <= r_data[26705];
                
                r_data[26707] <= r_data[26706];
                
                r_data[26708] <= r_data[26707];
                
                r_data[26709] <= r_data[26708];
                
                r_data[26710] <= r_data[26709];
                
                r_data[26711] <= r_data[26710];
                
                r_data[26712] <= r_data[26711];
                
                r_data[26713] <= r_data[26712];
                
                r_data[26714] <= r_data[26713];
                
                r_data[26715] <= r_data[26714];
                
                r_data[26716] <= r_data[26715];
                
                r_data[26717] <= r_data[26716];
                
                r_data[26718] <= r_data[26717];
                
                r_data[26719] <= r_data[26718];
                
                r_data[26720] <= r_data[26719];
                
                r_data[26721] <= r_data[26720];
                
                r_data[26722] <= r_data[26721];
                
                r_data[26723] <= r_data[26722];
                
                r_data[26724] <= r_data[26723];
                
                r_data[26725] <= r_data[26724];
                
                r_data[26726] <= r_data[26725];
                
                r_data[26727] <= r_data[26726];
                
                r_data[26728] <= r_data[26727];
                
                r_data[26729] <= r_data[26728];
                
                r_data[26730] <= r_data[26729];
                
                r_data[26731] <= r_data[26730];
                
                r_data[26732] <= r_data[26731];
                
                r_data[26733] <= r_data[26732];
                
                r_data[26734] <= r_data[26733];
                
                r_data[26735] <= r_data[26734];
                
                r_data[26736] <= r_data[26735];
                
                r_data[26737] <= r_data[26736];
                
                r_data[26738] <= r_data[26737];
                
                r_data[26739] <= r_data[26738];
                
                r_data[26740] <= r_data[26739];
                
                r_data[26741] <= r_data[26740];
                
                r_data[26742] <= r_data[26741];
                
                r_data[26743] <= r_data[26742];
                
                r_data[26744] <= r_data[26743];
                
                r_data[26745] <= r_data[26744];
                
                r_data[26746] <= r_data[26745];
                
                r_data[26747] <= r_data[26746];
                
                r_data[26748] <= r_data[26747];
                
                r_data[26749] <= r_data[26748];
                
                r_data[26750] <= r_data[26749];
                
                r_data[26751] <= r_data[26750];
                
                r_data[26752] <= r_data[26751];
                
                r_data[26753] <= r_data[26752];
                
                r_data[26754] <= r_data[26753];
                
                r_data[26755] <= r_data[26754];
                
                r_data[26756] <= r_data[26755];
                
                r_data[26757] <= r_data[26756];
                
                r_data[26758] <= r_data[26757];
                
                r_data[26759] <= r_data[26758];
                
                r_data[26760] <= r_data[26759];
                
                r_data[26761] <= r_data[26760];
                
                r_data[26762] <= r_data[26761];
                
                r_data[26763] <= r_data[26762];
                
                r_data[26764] <= r_data[26763];
                
                r_data[26765] <= r_data[26764];
                
                r_data[26766] <= r_data[26765];
                
                r_data[26767] <= r_data[26766];
                
                r_data[26768] <= r_data[26767];
                
                r_data[26769] <= r_data[26768];
                
                r_data[26770] <= r_data[26769];
                
                r_data[26771] <= r_data[26770];
                
                r_data[26772] <= r_data[26771];
                
                r_data[26773] <= r_data[26772];
                
                r_data[26774] <= r_data[26773];
                
                r_data[26775] <= r_data[26774];
                
                r_data[26776] <= r_data[26775];
                
                r_data[26777] <= r_data[26776];
                
                r_data[26778] <= r_data[26777];
                
                r_data[26779] <= r_data[26778];
                
                r_data[26780] <= r_data[26779];
                
                r_data[26781] <= r_data[26780];
                
                r_data[26782] <= r_data[26781];
                
                r_data[26783] <= r_data[26782];
                
                r_data[26784] <= r_data[26783];
                
                r_data[26785] <= r_data[26784];
                
                r_data[26786] <= r_data[26785];
                
                r_data[26787] <= r_data[26786];
                
                r_data[26788] <= r_data[26787];
                
                r_data[26789] <= r_data[26788];
                
                r_data[26790] <= r_data[26789];
                
                r_data[26791] <= r_data[26790];
                
                r_data[26792] <= r_data[26791];
                
                r_data[26793] <= r_data[26792];
                
                r_data[26794] <= r_data[26793];
                
                r_data[26795] <= r_data[26794];
                
                r_data[26796] <= r_data[26795];
                
                r_data[26797] <= r_data[26796];
                
                r_data[26798] <= r_data[26797];
                
                r_data[26799] <= r_data[26798];
                
                r_data[26800] <= r_data[26799];
                
                r_data[26801] <= r_data[26800];
                
                r_data[26802] <= r_data[26801];
                
                r_data[26803] <= r_data[26802];
                
                r_data[26804] <= r_data[26803];
                
                r_data[26805] <= r_data[26804];
                
                r_data[26806] <= r_data[26805];
                
                r_data[26807] <= r_data[26806];
                
                r_data[26808] <= r_data[26807];
                
                r_data[26809] <= r_data[26808];
                
                r_data[26810] <= r_data[26809];
                
                r_data[26811] <= r_data[26810];
                
                r_data[26812] <= r_data[26811];
                
                r_data[26813] <= r_data[26812];
                
                r_data[26814] <= r_data[26813];
                
                r_data[26815] <= r_data[26814];
                
                r_data[26816] <= r_data[26815];
                
                r_data[26817] <= r_data[26816];
                
                r_data[26818] <= r_data[26817];
                
                r_data[26819] <= r_data[26818];
                
                r_data[26820] <= r_data[26819];
                
                r_data[26821] <= r_data[26820];
                
                r_data[26822] <= r_data[26821];
                
                r_data[26823] <= r_data[26822];
                
                r_data[26824] <= r_data[26823];
                
                r_data[26825] <= r_data[26824];
                
                r_data[26826] <= r_data[26825];
                
                r_data[26827] <= r_data[26826];
                
                r_data[26828] <= r_data[26827];
                
                r_data[26829] <= r_data[26828];
                
                r_data[26830] <= r_data[26829];
                
                r_data[26831] <= r_data[26830];
                
                r_data[26832] <= r_data[26831];
                
                r_data[26833] <= r_data[26832];
                
                r_data[26834] <= r_data[26833];
                
                r_data[26835] <= r_data[26834];
                
                r_data[26836] <= r_data[26835];
                
                r_data[26837] <= r_data[26836];
                
                r_data[26838] <= r_data[26837];
                
                r_data[26839] <= r_data[26838];
                
                r_data[26840] <= r_data[26839];
                
                r_data[26841] <= r_data[26840];
                
                r_data[26842] <= r_data[26841];
                
                r_data[26843] <= r_data[26842];
                
                r_data[26844] <= r_data[26843];
                
                r_data[26845] <= r_data[26844];
                
                r_data[26846] <= r_data[26845];
                
                r_data[26847] <= r_data[26846];
                
                r_data[26848] <= r_data[26847];
                
                r_data[26849] <= r_data[26848];
                
                r_data[26850] <= r_data[26849];
                
                r_data[26851] <= r_data[26850];
                
                r_data[26852] <= r_data[26851];
                
                r_data[26853] <= r_data[26852];
                
                r_data[26854] <= r_data[26853];
                
                r_data[26855] <= r_data[26854];
                
                r_data[26856] <= r_data[26855];
                
                r_data[26857] <= r_data[26856];
                
                r_data[26858] <= r_data[26857];
                
                r_data[26859] <= r_data[26858];
                
                r_data[26860] <= r_data[26859];
                
                r_data[26861] <= r_data[26860];
                
                r_data[26862] <= r_data[26861];
                
                r_data[26863] <= r_data[26862];
                
                r_data[26864] <= r_data[26863];
                
                r_data[26865] <= r_data[26864];
                
                r_data[26866] <= r_data[26865];
                
                r_data[26867] <= r_data[26866];
                
                r_data[26868] <= r_data[26867];
                
                r_data[26869] <= r_data[26868];
                
                r_data[26870] <= r_data[26869];
                
                r_data[26871] <= r_data[26870];
                
                r_data[26872] <= r_data[26871];
                
                r_data[26873] <= r_data[26872];
                
                r_data[26874] <= r_data[26873];
                
                r_data[26875] <= r_data[26874];
                
                r_data[26876] <= r_data[26875];
                
                r_data[26877] <= r_data[26876];
                
                r_data[26878] <= r_data[26877];
                
                r_data[26879] <= r_data[26878];
                
                r_data[26880] <= r_data[26879];
                
                r_data[26881] <= r_data[26880];
                
                r_data[26882] <= r_data[26881];
                
                r_data[26883] <= r_data[26882];
                
                r_data[26884] <= r_data[26883];
                
                r_data[26885] <= r_data[26884];
                
                r_data[26886] <= r_data[26885];
                
                r_data[26887] <= r_data[26886];
                
                r_data[26888] <= r_data[26887];
                
                r_data[26889] <= r_data[26888];
                
                r_data[26890] <= r_data[26889];
                
                r_data[26891] <= r_data[26890];
                
                r_data[26892] <= r_data[26891];
                
                r_data[26893] <= r_data[26892];
                
                r_data[26894] <= r_data[26893];
                
                r_data[26895] <= r_data[26894];
                
                r_data[26896] <= r_data[26895];
                
                r_data[26897] <= r_data[26896];
                
                r_data[26898] <= r_data[26897];
                
                r_data[26899] <= r_data[26898];
                
                r_data[26900] <= r_data[26899];
                
                r_data[26901] <= r_data[26900];
                
                r_data[26902] <= r_data[26901];
                
                r_data[26903] <= r_data[26902];
                
                r_data[26904] <= r_data[26903];
                
                r_data[26905] <= r_data[26904];
                
                r_data[26906] <= r_data[26905];
                
                r_data[26907] <= r_data[26906];
                
                r_data[26908] <= r_data[26907];
                
                r_data[26909] <= r_data[26908];
                
                r_data[26910] <= r_data[26909];
                
                r_data[26911] <= r_data[26910];
                
                r_data[26912] <= r_data[26911];
                
                r_data[26913] <= r_data[26912];
                
                r_data[26914] <= r_data[26913];
                
                r_data[26915] <= r_data[26914];
                
                r_data[26916] <= r_data[26915];
                
                r_data[26917] <= r_data[26916];
                
                r_data[26918] <= r_data[26917];
                
                r_data[26919] <= r_data[26918];
                
                r_data[26920] <= r_data[26919];
                
                r_data[26921] <= r_data[26920];
                
                r_data[26922] <= r_data[26921];
                
                r_data[26923] <= r_data[26922];
                
                r_data[26924] <= r_data[26923];
                
                r_data[26925] <= r_data[26924];
                
                r_data[26926] <= r_data[26925];
                
                r_data[26927] <= r_data[26926];
                
                r_data[26928] <= r_data[26927];
                
                r_data[26929] <= r_data[26928];
                
                r_data[26930] <= r_data[26929];
                
                r_data[26931] <= r_data[26930];
                
                r_data[26932] <= r_data[26931];
                
                r_data[26933] <= r_data[26932];
                
                r_data[26934] <= r_data[26933];
                
                r_data[26935] <= r_data[26934];
                
                r_data[26936] <= r_data[26935];
                
                r_data[26937] <= r_data[26936];
                
                r_data[26938] <= r_data[26937];
                
                r_data[26939] <= r_data[26938];
                
                r_data[26940] <= r_data[26939];
                
                r_data[26941] <= r_data[26940];
                
                r_data[26942] <= r_data[26941];
                
                r_data[26943] <= r_data[26942];
                
                r_data[26944] <= r_data[26943];
                
                r_data[26945] <= r_data[26944];
                
                r_data[26946] <= r_data[26945];
                
                r_data[26947] <= r_data[26946];
                
                r_data[26948] <= r_data[26947];
                
                r_data[26949] <= r_data[26948];
                
                r_data[26950] <= r_data[26949];
                
                r_data[26951] <= r_data[26950];
                
                r_data[26952] <= r_data[26951];
                
                r_data[26953] <= r_data[26952];
                
                r_data[26954] <= r_data[26953];
                
                r_data[26955] <= r_data[26954];
                
                r_data[26956] <= r_data[26955];
                
                r_data[26957] <= r_data[26956];
                
                r_data[26958] <= r_data[26957];
                
                r_data[26959] <= r_data[26958];
                
                r_data[26960] <= r_data[26959];
                
                r_data[26961] <= r_data[26960];
                
                r_data[26962] <= r_data[26961];
                
                r_data[26963] <= r_data[26962];
                
                r_data[26964] <= r_data[26963];
                
                r_data[26965] <= r_data[26964];
                
                r_data[26966] <= r_data[26965];
                
                r_data[26967] <= r_data[26966];
                
                r_data[26968] <= r_data[26967];
                
                r_data[26969] <= r_data[26968];
                
                r_data[26970] <= r_data[26969];
                
                r_data[26971] <= r_data[26970];
                
                r_data[26972] <= r_data[26971];
                
                r_data[26973] <= r_data[26972];
                
                r_data[26974] <= r_data[26973];
                
                r_data[26975] <= r_data[26974];
                
                r_data[26976] <= r_data[26975];
                
                r_data[26977] <= r_data[26976];
                
                r_data[26978] <= r_data[26977];
                
                r_data[26979] <= r_data[26978];
                
                r_data[26980] <= r_data[26979];
                
                r_data[26981] <= r_data[26980];
                
                r_data[26982] <= r_data[26981];
                
                r_data[26983] <= r_data[26982];
                
                r_data[26984] <= r_data[26983];
                
                r_data[26985] <= r_data[26984];
                
                r_data[26986] <= r_data[26985];
                
                r_data[26987] <= r_data[26986];
                
                r_data[26988] <= r_data[26987];
                
                r_data[26989] <= r_data[26988];
                
                r_data[26990] <= r_data[26989];
                
                r_data[26991] <= r_data[26990];
                
                r_data[26992] <= r_data[26991];
                
                r_data[26993] <= r_data[26992];
                
                r_data[26994] <= r_data[26993];
                
                r_data[26995] <= r_data[26994];
                
                r_data[26996] <= r_data[26995];
                
                r_data[26997] <= r_data[26996];
                
                r_data[26998] <= r_data[26997];
                
                r_data[26999] <= r_data[26998];
                
                r_data[27000] <= r_data[26999];
                
                r_data[27001] <= r_data[27000];
                
                r_data[27002] <= r_data[27001];
                
                r_data[27003] <= r_data[27002];
                
                r_data[27004] <= r_data[27003];
                
                r_data[27005] <= r_data[27004];
                
                r_data[27006] <= r_data[27005];
                
                r_data[27007] <= r_data[27006];
                
                r_data[27008] <= r_data[27007];
                
                r_data[27009] <= r_data[27008];
                
                r_data[27010] <= r_data[27009];
                
                r_data[27011] <= r_data[27010];
                
                r_data[27012] <= r_data[27011];
                
                r_data[27013] <= r_data[27012];
                
                r_data[27014] <= r_data[27013];
                
                r_data[27015] <= r_data[27014];
                
                r_data[27016] <= r_data[27015];
                
                r_data[27017] <= r_data[27016];
                
                r_data[27018] <= r_data[27017];
                
                r_data[27019] <= r_data[27018];
                
                r_data[27020] <= r_data[27019];
                
                r_data[27021] <= r_data[27020];
                
                r_data[27022] <= r_data[27021];
                
                r_data[27023] <= r_data[27022];
                
                r_data[27024] <= r_data[27023];
                
                r_data[27025] <= r_data[27024];
                
                r_data[27026] <= r_data[27025];
                
                r_data[27027] <= r_data[27026];
                
                r_data[27028] <= r_data[27027];
                
                r_data[27029] <= r_data[27028];
                
                r_data[27030] <= r_data[27029];
                
                r_data[27031] <= r_data[27030];
                
                r_data[27032] <= r_data[27031];
                
                r_data[27033] <= r_data[27032];
                
                r_data[27034] <= r_data[27033];
                
                r_data[27035] <= r_data[27034];
                
                r_data[27036] <= r_data[27035];
                
                r_data[27037] <= r_data[27036];
                
                r_data[27038] <= r_data[27037];
                
                r_data[27039] <= r_data[27038];
                
                r_data[27040] <= r_data[27039];
                
                r_data[27041] <= r_data[27040];
                
                r_data[27042] <= r_data[27041];
                
                r_data[27043] <= r_data[27042];
                
                r_data[27044] <= r_data[27043];
                
                r_data[27045] <= r_data[27044];
                
                r_data[27046] <= r_data[27045];
                
                r_data[27047] <= r_data[27046];
                
                r_data[27048] <= r_data[27047];
                
                r_data[27049] <= r_data[27048];
                
                r_data[27050] <= r_data[27049];
                
                r_data[27051] <= r_data[27050];
                
                r_data[27052] <= r_data[27051];
                
                r_data[27053] <= r_data[27052];
                
                r_data[27054] <= r_data[27053];
                
                r_data[27055] <= r_data[27054];
                
                r_data[27056] <= r_data[27055];
                
                r_data[27057] <= r_data[27056];
                
                r_data[27058] <= r_data[27057];
                
                r_data[27059] <= r_data[27058];
                
                r_data[27060] <= r_data[27059];
                
                r_data[27061] <= r_data[27060];
                
                r_data[27062] <= r_data[27061];
                
                r_data[27063] <= r_data[27062];
                
                r_data[27064] <= r_data[27063];
                
                r_data[27065] <= r_data[27064];
                
                r_data[27066] <= r_data[27065];
                
                r_data[27067] <= r_data[27066];
                
                r_data[27068] <= r_data[27067];
                
                r_data[27069] <= r_data[27068];
                
                r_data[27070] <= r_data[27069];
                
                r_data[27071] <= r_data[27070];
                
                r_data[27072] <= r_data[27071];
                
                r_data[27073] <= r_data[27072];
                
                r_data[27074] <= r_data[27073];
                
                r_data[27075] <= r_data[27074];
                
                r_data[27076] <= r_data[27075];
                
                r_data[27077] <= r_data[27076];
                
                r_data[27078] <= r_data[27077];
                
                r_data[27079] <= r_data[27078];
                
                r_data[27080] <= r_data[27079];
                
                r_data[27081] <= r_data[27080];
                
                r_data[27082] <= r_data[27081];
                
                r_data[27083] <= r_data[27082];
                
                r_data[27084] <= r_data[27083];
                
                r_data[27085] <= r_data[27084];
                
                r_data[27086] <= r_data[27085];
                
                r_data[27087] <= r_data[27086];
                
                r_data[27088] <= r_data[27087];
                
                r_data[27089] <= r_data[27088];
                
                r_data[27090] <= r_data[27089];
                
                r_data[27091] <= r_data[27090];
                
                r_data[27092] <= r_data[27091];
                
                r_data[27093] <= r_data[27092];
                
                r_data[27094] <= r_data[27093];
                
                r_data[27095] <= r_data[27094];
                
                r_data[27096] <= r_data[27095];
                
                r_data[27097] <= r_data[27096];
                
                r_data[27098] <= r_data[27097];
                
                r_data[27099] <= r_data[27098];
                
                r_data[27100] <= r_data[27099];
                
                r_data[27101] <= r_data[27100];
                
                r_data[27102] <= r_data[27101];
                
                r_data[27103] <= r_data[27102];
                
                r_data[27104] <= r_data[27103];
                
                r_data[27105] <= r_data[27104];
                
                r_data[27106] <= r_data[27105];
                
                r_data[27107] <= r_data[27106];
                
                r_data[27108] <= r_data[27107];
                
                r_data[27109] <= r_data[27108];
                
                r_data[27110] <= r_data[27109];
                
                r_data[27111] <= r_data[27110];
                
                r_data[27112] <= r_data[27111];
                
                r_data[27113] <= r_data[27112];
                
                r_data[27114] <= r_data[27113];
                
                r_data[27115] <= r_data[27114];
                
                r_data[27116] <= r_data[27115];
                
                r_data[27117] <= r_data[27116];
                
                r_data[27118] <= r_data[27117];
                
                r_data[27119] <= r_data[27118];
                
                r_data[27120] <= r_data[27119];
                
                r_data[27121] <= r_data[27120];
                
                r_data[27122] <= r_data[27121];
                
                r_data[27123] <= r_data[27122];
                
                r_data[27124] <= r_data[27123];
                
                r_data[27125] <= r_data[27124];
                
                r_data[27126] <= r_data[27125];
                
                r_data[27127] <= r_data[27126];
                
                r_data[27128] <= r_data[27127];
                
                r_data[27129] <= r_data[27128];
                
                r_data[27130] <= r_data[27129];
                
                r_data[27131] <= r_data[27130];
                
                r_data[27132] <= r_data[27131];
                
                r_data[27133] <= r_data[27132];
                
                r_data[27134] <= r_data[27133];
                
                r_data[27135] <= r_data[27134];
                
                r_data[27136] <= r_data[27135];
                
                r_data[27137] <= r_data[27136];
                
                r_data[27138] <= r_data[27137];
                
                r_data[27139] <= r_data[27138];
                
                r_data[27140] <= r_data[27139];
                
                r_data[27141] <= r_data[27140];
                
                r_data[27142] <= r_data[27141];
                
                r_data[27143] <= r_data[27142];
                
                r_data[27144] <= r_data[27143];
                
                r_data[27145] <= r_data[27144];
                
                r_data[27146] <= r_data[27145];
                
                r_data[27147] <= r_data[27146];
                
                r_data[27148] <= r_data[27147];
                
                r_data[27149] <= r_data[27148];
                
                r_data[27150] <= r_data[27149];
                
                r_data[27151] <= r_data[27150];
                
                r_data[27152] <= r_data[27151];
                
                r_data[27153] <= r_data[27152];
                
                r_data[27154] <= r_data[27153];
                
                r_data[27155] <= r_data[27154];
                
                r_data[27156] <= r_data[27155];
                
                r_data[27157] <= r_data[27156];
                
                r_data[27158] <= r_data[27157];
                
                r_data[27159] <= r_data[27158];
                
                r_data[27160] <= r_data[27159];
                
                r_data[27161] <= r_data[27160];
                
                r_data[27162] <= r_data[27161];
                
                r_data[27163] <= r_data[27162];
                
                r_data[27164] <= r_data[27163];
                
                r_data[27165] <= r_data[27164];
                
                r_data[27166] <= r_data[27165];
                
                r_data[27167] <= r_data[27166];
                
                r_data[27168] <= r_data[27167];
                
                r_data[27169] <= r_data[27168];
                
                r_data[27170] <= r_data[27169];
                
                r_data[27171] <= r_data[27170];
                
                r_data[27172] <= r_data[27171];
                
                r_data[27173] <= r_data[27172];
                
                r_data[27174] <= r_data[27173];
                
                r_data[27175] <= r_data[27174];
                
                r_data[27176] <= r_data[27175];
                
                r_data[27177] <= r_data[27176];
                
                r_data[27178] <= r_data[27177];
                
                r_data[27179] <= r_data[27178];
                
                r_data[27180] <= r_data[27179];
                
                r_data[27181] <= r_data[27180];
                
                r_data[27182] <= r_data[27181];
                
                r_data[27183] <= r_data[27182];
                
                r_data[27184] <= r_data[27183];
                
                r_data[27185] <= r_data[27184];
                
                r_data[27186] <= r_data[27185];
                
                r_data[27187] <= r_data[27186];
                
                r_data[27188] <= r_data[27187];
                
                r_data[27189] <= r_data[27188];
                
                r_data[27190] <= r_data[27189];
                
                r_data[27191] <= r_data[27190];
                
                r_data[27192] <= r_data[27191];
                
                r_data[27193] <= r_data[27192];
                
                r_data[27194] <= r_data[27193];
                
                r_data[27195] <= r_data[27194];
                
                r_data[27196] <= r_data[27195];
                
                r_data[27197] <= r_data[27196];
                
                r_data[27198] <= r_data[27197];
                
                r_data[27199] <= r_data[27198];
                
                r_data[27200] <= r_data[27199];
                
                r_data[27201] <= r_data[27200];
                
                r_data[27202] <= r_data[27201];
                
                r_data[27203] <= r_data[27202];
                
                r_data[27204] <= r_data[27203];
                
                r_data[27205] <= r_data[27204];
                
                r_data[27206] <= r_data[27205];
                
                r_data[27207] <= r_data[27206];
                
                r_data[27208] <= r_data[27207];
                
                r_data[27209] <= r_data[27208];
                
                r_data[27210] <= r_data[27209];
                
                r_data[27211] <= r_data[27210];
                
                r_data[27212] <= r_data[27211];
                
                r_data[27213] <= r_data[27212];
                
                r_data[27214] <= r_data[27213];
                
                r_data[27215] <= r_data[27214];
                
                r_data[27216] <= r_data[27215];
                
                r_data[27217] <= r_data[27216];
                
                r_data[27218] <= r_data[27217];
                
                r_data[27219] <= r_data[27218];
                
                r_data[27220] <= r_data[27219];
                
                r_data[27221] <= r_data[27220];
                
                r_data[27222] <= r_data[27221];
                
                r_data[27223] <= r_data[27222];
                
                r_data[27224] <= r_data[27223];
                
                r_data[27225] <= r_data[27224];
                
                r_data[27226] <= r_data[27225];
                
                r_data[27227] <= r_data[27226];
                
                r_data[27228] <= r_data[27227];
                
                r_data[27229] <= r_data[27228];
                
                r_data[27230] <= r_data[27229];
                
                r_data[27231] <= r_data[27230];
                
                r_data[27232] <= r_data[27231];
                
                r_data[27233] <= r_data[27232];
                
                r_data[27234] <= r_data[27233];
                
                r_data[27235] <= r_data[27234];
                
                r_data[27236] <= r_data[27235];
                
                r_data[27237] <= r_data[27236];
                
                r_data[27238] <= r_data[27237];
                
                r_data[27239] <= r_data[27238];
                
                r_data[27240] <= r_data[27239];
                
                r_data[27241] <= r_data[27240];
                
                r_data[27242] <= r_data[27241];
                
                r_data[27243] <= r_data[27242];
                
                r_data[27244] <= r_data[27243];
                
                r_data[27245] <= r_data[27244];
                
                r_data[27246] <= r_data[27245];
                
                r_data[27247] <= r_data[27246];
                
                r_data[27248] <= r_data[27247];
                
                r_data[27249] <= r_data[27248];
                
                r_data[27250] <= r_data[27249];
                
                r_data[27251] <= r_data[27250];
                
                r_data[27252] <= r_data[27251];
                
                r_data[27253] <= r_data[27252];
                
                r_data[27254] <= r_data[27253];
                
                r_data[27255] <= r_data[27254];
                
                r_data[27256] <= r_data[27255];
                
                r_data[27257] <= r_data[27256];
                
                r_data[27258] <= r_data[27257];
                
                r_data[27259] <= r_data[27258];
                
                r_data[27260] <= r_data[27259];
                
                r_data[27261] <= r_data[27260];
                
                r_data[27262] <= r_data[27261];
                
                r_data[27263] <= r_data[27262];
                
                r_data[27264] <= r_data[27263];
                
                r_data[27265] <= r_data[27264];
                
                r_data[27266] <= r_data[27265];
                
                r_data[27267] <= r_data[27266];
                
                r_data[27268] <= r_data[27267];
                
                r_data[27269] <= r_data[27268];
                
                r_data[27270] <= r_data[27269];
                
                r_data[27271] <= r_data[27270];
                
                r_data[27272] <= r_data[27271];
                
                r_data[27273] <= r_data[27272];
                
                r_data[27274] <= r_data[27273];
                
                r_data[27275] <= r_data[27274];
                
                r_data[27276] <= r_data[27275];
                
                r_data[27277] <= r_data[27276];
                
                r_data[27278] <= r_data[27277];
                
                r_data[27279] <= r_data[27278];
                
                r_data[27280] <= r_data[27279];
                
                r_data[27281] <= r_data[27280];
                
                r_data[27282] <= r_data[27281];
                
                r_data[27283] <= r_data[27282];
                
                r_data[27284] <= r_data[27283];
                
                r_data[27285] <= r_data[27284];
                
                r_data[27286] <= r_data[27285];
                
                r_data[27287] <= r_data[27286];
                
                r_data[27288] <= r_data[27287];
                
                r_data[27289] <= r_data[27288];
                
                r_data[27290] <= r_data[27289];
                
                r_data[27291] <= r_data[27290];
                
                r_data[27292] <= r_data[27291];
                
                r_data[27293] <= r_data[27292];
                
                r_data[27294] <= r_data[27293];
                
                r_data[27295] <= r_data[27294];
                
                r_data[27296] <= r_data[27295];
                
                r_data[27297] <= r_data[27296];
                
                r_data[27298] <= r_data[27297];
                
                r_data[27299] <= r_data[27298];
                
                r_data[27300] <= r_data[27299];
                
                r_data[27301] <= r_data[27300];
                
                r_data[27302] <= r_data[27301];
                
                r_data[27303] <= r_data[27302];
                
                r_data[27304] <= r_data[27303];
                
                r_data[27305] <= r_data[27304];
                
                r_data[27306] <= r_data[27305];
                
                r_data[27307] <= r_data[27306];
                
                r_data[27308] <= r_data[27307];
                
                r_data[27309] <= r_data[27308];
                
                r_data[27310] <= r_data[27309];
                
                r_data[27311] <= r_data[27310];
                
                r_data[27312] <= r_data[27311];
                
                r_data[27313] <= r_data[27312];
                
                r_data[27314] <= r_data[27313];
                
                r_data[27315] <= r_data[27314];
                
                r_data[27316] <= r_data[27315];
                
                r_data[27317] <= r_data[27316];
                
                r_data[27318] <= r_data[27317];
                
                r_data[27319] <= r_data[27318];
                
                r_data[27320] <= r_data[27319];
                
                r_data[27321] <= r_data[27320];
                
                r_data[27322] <= r_data[27321];
                
                r_data[27323] <= r_data[27322];
                
                r_data[27324] <= r_data[27323];
                
                r_data[27325] <= r_data[27324];
                
                r_data[27326] <= r_data[27325];
                
                r_data[27327] <= r_data[27326];
                
                r_data[27328] <= r_data[27327];
                
                r_data[27329] <= r_data[27328];
                
                r_data[27330] <= r_data[27329];
                
                r_data[27331] <= r_data[27330];
                
                r_data[27332] <= r_data[27331];
                
                r_data[27333] <= r_data[27332];
                
                r_data[27334] <= r_data[27333];
                
                r_data[27335] <= r_data[27334];
                
                r_data[27336] <= r_data[27335];
                
                r_data[27337] <= r_data[27336];
                
                r_data[27338] <= r_data[27337];
                
                r_data[27339] <= r_data[27338];
                
                r_data[27340] <= r_data[27339];
                
                r_data[27341] <= r_data[27340];
                
                r_data[27342] <= r_data[27341];
                
                r_data[27343] <= r_data[27342];
                
                r_data[27344] <= r_data[27343];
                
                r_data[27345] <= r_data[27344];
                
                r_data[27346] <= r_data[27345];
                
                r_data[27347] <= r_data[27346];
                
                r_data[27348] <= r_data[27347];
                
                r_data[27349] <= r_data[27348];
                
                r_data[27350] <= r_data[27349];
                
                r_data[27351] <= r_data[27350];
                
                r_data[27352] <= r_data[27351];
                
                r_data[27353] <= r_data[27352];
                
                r_data[27354] <= r_data[27353];
                
                r_data[27355] <= r_data[27354];
                
                r_data[27356] <= r_data[27355];
                
                r_data[27357] <= r_data[27356];
                
                r_data[27358] <= r_data[27357];
                
                r_data[27359] <= r_data[27358];
                
                r_data[27360] <= r_data[27359];
                
                r_data[27361] <= r_data[27360];
                
                r_data[27362] <= r_data[27361];
                
                r_data[27363] <= r_data[27362];
                
                r_data[27364] <= r_data[27363];
                
                r_data[27365] <= r_data[27364];
                
                r_data[27366] <= r_data[27365];
                
                r_data[27367] <= r_data[27366];
                
                r_data[27368] <= r_data[27367];
                
                r_data[27369] <= r_data[27368];
                
                r_data[27370] <= r_data[27369];
                
                r_data[27371] <= r_data[27370];
                
                r_data[27372] <= r_data[27371];
                
                r_data[27373] <= r_data[27372];
                
                r_data[27374] <= r_data[27373];
                
                r_data[27375] <= r_data[27374];
                
                r_data[27376] <= r_data[27375];
                
                r_data[27377] <= r_data[27376];
                
                r_data[27378] <= r_data[27377];
                
                r_data[27379] <= r_data[27378];
                
                r_data[27380] <= r_data[27379];
                
                r_data[27381] <= r_data[27380];
                
                r_data[27382] <= r_data[27381];
                
                r_data[27383] <= r_data[27382];
                
                r_data[27384] <= r_data[27383];
                
                r_data[27385] <= r_data[27384];
                
                r_data[27386] <= r_data[27385];
                
                r_data[27387] <= r_data[27386];
                
                r_data[27388] <= r_data[27387];
                
                r_data[27389] <= r_data[27388];
                
                r_data[27390] <= r_data[27389];
                
                r_data[27391] <= r_data[27390];
                
                r_data[27392] <= r_data[27391];
                
                r_data[27393] <= r_data[27392];
                
                r_data[27394] <= r_data[27393];
                
                r_data[27395] <= r_data[27394];
                
                r_data[27396] <= r_data[27395];
                
                r_data[27397] <= r_data[27396];
                
                r_data[27398] <= r_data[27397];
                
                r_data[27399] <= r_data[27398];
                
                r_data[27400] <= r_data[27399];
                
                r_data[27401] <= r_data[27400];
                
                r_data[27402] <= r_data[27401];
                
                r_data[27403] <= r_data[27402];
                
                r_data[27404] <= r_data[27403];
                
                r_data[27405] <= r_data[27404];
                
                r_data[27406] <= r_data[27405];
                
                r_data[27407] <= r_data[27406];
                
                r_data[27408] <= r_data[27407];
                
                r_data[27409] <= r_data[27408];
                
                r_data[27410] <= r_data[27409];
                
                r_data[27411] <= r_data[27410];
                
                r_data[27412] <= r_data[27411];
                
                r_data[27413] <= r_data[27412];
                
                r_data[27414] <= r_data[27413];
                
                r_data[27415] <= r_data[27414];
                
                r_data[27416] <= r_data[27415];
                
                r_data[27417] <= r_data[27416];
                
                r_data[27418] <= r_data[27417];
                
                r_data[27419] <= r_data[27418];
                
                r_data[27420] <= r_data[27419];
                
                r_data[27421] <= r_data[27420];
                
                r_data[27422] <= r_data[27421];
                
                r_data[27423] <= r_data[27422];
                
                r_data[27424] <= r_data[27423];
                
                r_data[27425] <= r_data[27424];
                
                r_data[27426] <= r_data[27425];
                
                r_data[27427] <= r_data[27426];
                
                r_data[27428] <= r_data[27427];
                
                r_data[27429] <= r_data[27428];
                
                r_data[27430] <= r_data[27429];
                
                r_data[27431] <= r_data[27430];
                
                r_data[27432] <= r_data[27431];
                
                r_data[27433] <= r_data[27432];
                
                r_data[27434] <= r_data[27433];
                
                r_data[27435] <= r_data[27434];
                
                r_data[27436] <= r_data[27435];
                
                r_data[27437] <= r_data[27436];
                
                r_data[27438] <= r_data[27437];
                
                r_data[27439] <= r_data[27438];
                
                r_data[27440] <= r_data[27439];
                
                r_data[27441] <= r_data[27440];
                
                r_data[27442] <= r_data[27441];
                
                r_data[27443] <= r_data[27442];
                
                r_data[27444] <= r_data[27443];
                
                r_data[27445] <= r_data[27444];
                
                r_data[27446] <= r_data[27445];
                
                r_data[27447] <= r_data[27446];
                
                r_data[27448] <= r_data[27447];
                
                r_data[27449] <= r_data[27448];
                
                r_data[27450] <= r_data[27449];
                
                r_data[27451] <= r_data[27450];
                
                r_data[27452] <= r_data[27451];
                
                r_data[27453] <= r_data[27452];
                
                r_data[27454] <= r_data[27453];
                
                r_data[27455] <= r_data[27454];
                
                r_data[27456] <= r_data[27455];
                
                r_data[27457] <= r_data[27456];
                
                r_data[27458] <= r_data[27457];
                
                r_data[27459] <= r_data[27458];
                
                r_data[27460] <= r_data[27459];
                
                r_data[27461] <= r_data[27460];
                
                r_data[27462] <= r_data[27461];
                
                r_data[27463] <= r_data[27462];
                
                r_data[27464] <= r_data[27463];
                
                r_data[27465] <= r_data[27464];
                
                r_data[27466] <= r_data[27465];
                
                r_data[27467] <= r_data[27466];
                
                r_data[27468] <= r_data[27467];
                
                r_data[27469] <= r_data[27468];
                
                r_data[27470] <= r_data[27469];
                
                r_data[27471] <= r_data[27470];
                
                r_data[27472] <= r_data[27471];
                
                r_data[27473] <= r_data[27472];
                
                r_data[27474] <= r_data[27473];
                
                r_data[27475] <= r_data[27474];
                
                r_data[27476] <= r_data[27475];
                
                r_data[27477] <= r_data[27476];
                
                r_data[27478] <= r_data[27477];
                
                r_data[27479] <= r_data[27478];
                
                r_data[27480] <= r_data[27479];
                
                r_data[27481] <= r_data[27480];
                
                r_data[27482] <= r_data[27481];
                
                r_data[27483] <= r_data[27482];
                
                r_data[27484] <= r_data[27483];
                
                r_data[27485] <= r_data[27484];
                
                r_data[27486] <= r_data[27485];
                
                r_data[27487] <= r_data[27486];
                
                r_data[27488] <= r_data[27487];
                
                r_data[27489] <= r_data[27488];
                
                r_data[27490] <= r_data[27489];
                
                r_data[27491] <= r_data[27490];
                
                r_data[27492] <= r_data[27491];
                
                r_data[27493] <= r_data[27492];
                
                r_data[27494] <= r_data[27493];
                
                r_data[27495] <= r_data[27494];
                
                r_data[27496] <= r_data[27495];
                
                r_data[27497] <= r_data[27496];
                
                r_data[27498] <= r_data[27497];
                
                r_data[27499] <= r_data[27498];
                
                r_data[27500] <= r_data[27499];
                
                r_data[27501] <= r_data[27500];
                
                r_data[27502] <= r_data[27501];
                
                r_data[27503] <= r_data[27502];
                
                r_data[27504] <= r_data[27503];
                
                r_data[27505] <= r_data[27504];
                
                r_data[27506] <= r_data[27505];
                
                r_data[27507] <= r_data[27506];
                
                r_data[27508] <= r_data[27507];
                
                r_data[27509] <= r_data[27508];
                
                r_data[27510] <= r_data[27509];
                
                r_data[27511] <= r_data[27510];
                
                r_data[27512] <= r_data[27511];
                
                r_data[27513] <= r_data[27512];
                
                r_data[27514] <= r_data[27513];
                
                r_data[27515] <= r_data[27514];
                
                r_data[27516] <= r_data[27515];
                
                r_data[27517] <= r_data[27516];
                
                r_data[27518] <= r_data[27517];
                
                r_data[27519] <= r_data[27518];
                
                r_data[27520] <= r_data[27519];
                
                r_data[27521] <= r_data[27520];
                
                r_data[27522] <= r_data[27521];
                
                r_data[27523] <= r_data[27522];
                
                r_data[27524] <= r_data[27523];
                
                r_data[27525] <= r_data[27524];
                
                r_data[27526] <= r_data[27525];
                
                r_data[27527] <= r_data[27526];
                
                r_data[27528] <= r_data[27527];
                
                r_data[27529] <= r_data[27528];
                
                r_data[27530] <= r_data[27529];
                
                r_data[27531] <= r_data[27530];
                
                r_data[27532] <= r_data[27531];
                
                r_data[27533] <= r_data[27532];
                
                r_data[27534] <= r_data[27533];
                
                r_data[27535] <= r_data[27534];
                
                r_data[27536] <= r_data[27535];
                
                r_data[27537] <= r_data[27536];
                
                r_data[27538] <= r_data[27537];
                
                r_data[27539] <= r_data[27538];
                
                r_data[27540] <= r_data[27539];
                
                r_data[27541] <= r_data[27540];
                
                r_data[27542] <= r_data[27541];
                
                r_data[27543] <= r_data[27542];
                
                r_data[27544] <= r_data[27543];
                
                r_data[27545] <= r_data[27544];
                
                r_data[27546] <= r_data[27545];
                
                r_data[27547] <= r_data[27546];
                
                r_data[27548] <= r_data[27547];
                
                r_data[27549] <= r_data[27548];
                
                r_data[27550] <= r_data[27549];
                
                r_data[27551] <= r_data[27550];
                
                r_data[27552] <= r_data[27551];
                
                r_data[27553] <= r_data[27552];
                
                r_data[27554] <= r_data[27553];
                
                r_data[27555] <= r_data[27554];
                
                r_data[27556] <= r_data[27555];
                
                r_data[27557] <= r_data[27556];
                
                r_data[27558] <= r_data[27557];
                
                r_data[27559] <= r_data[27558];
                
                r_data[27560] <= r_data[27559];
                
                r_data[27561] <= r_data[27560];
                
                r_data[27562] <= r_data[27561];
                
                r_data[27563] <= r_data[27562];
                
                r_data[27564] <= r_data[27563];
                
                r_data[27565] <= r_data[27564];
                
                r_data[27566] <= r_data[27565];
                
                r_data[27567] <= r_data[27566];
                
                r_data[27568] <= r_data[27567];
                
                r_data[27569] <= r_data[27568];
                
                r_data[27570] <= r_data[27569];
                
                r_data[27571] <= r_data[27570];
                
                r_data[27572] <= r_data[27571];
                
                r_data[27573] <= r_data[27572];
                
                r_data[27574] <= r_data[27573];
                
                r_data[27575] <= r_data[27574];
                
                r_data[27576] <= r_data[27575];
                
                r_data[27577] <= r_data[27576];
                
                r_data[27578] <= r_data[27577];
                
                r_data[27579] <= r_data[27578];
                
                r_data[27580] <= r_data[27579];
                
                r_data[27581] <= r_data[27580];
                
                r_data[27582] <= r_data[27581];
                
                r_data[27583] <= r_data[27582];
                
                r_data[27584] <= r_data[27583];
                
                r_data[27585] <= r_data[27584];
                
                r_data[27586] <= r_data[27585];
                
                r_data[27587] <= r_data[27586];
                
                r_data[27588] <= r_data[27587];
                
                r_data[27589] <= r_data[27588];
                
                r_data[27590] <= r_data[27589];
                
                r_data[27591] <= r_data[27590];
                
                r_data[27592] <= r_data[27591];
                
                r_data[27593] <= r_data[27592];
                
                r_data[27594] <= r_data[27593];
                
                r_data[27595] <= r_data[27594];
                
                r_data[27596] <= r_data[27595];
                
                r_data[27597] <= r_data[27596];
                
                r_data[27598] <= r_data[27597];
                
                r_data[27599] <= r_data[27598];
                
                r_data[27600] <= r_data[27599];
                
                r_data[27601] <= r_data[27600];
                
                r_data[27602] <= r_data[27601];
                
                r_data[27603] <= r_data[27602];
                
                r_data[27604] <= r_data[27603];
                
                r_data[27605] <= r_data[27604];
                
                r_data[27606] <= r_data[27605];
                
                r_data[27607] <= r_data[27606];
                
                r_data[27608] <= r_data[27607];
                
                r_data[27609] <= r_data[27608];
                
                r_data[27610] <= r_data[27609];
                
                r_data[27611] <= r_data[27610];
                
                r_data[27612] <= r_data[27611];
                
                r_data[27613] <= r_data[27612];
                
                r_data[27614] <= r_data[27613];
                
                r_data[27615] <= r_data[27614];
                
                r_data[27616] <= r_data[27615];
                
                r_data[27617] <= r_data[27616];
                
                r_data[27618] <= r_data[27617];
                
                r_data[27619] <= r_data[27618];
                
                r_data[27620] <= r_data[27619];
                
                r_data[27621] <= r_data[27620];
                
                r_data[27622] <= r_data[27621];
                
                r_data[27623] <= r_data[27622];
                
                r_data[27624] <= r_data[27623];
                
                r_data[27625] <= r_data[27624];
                
                r_data[27626] <= r_data[27625];
                
                r_data[27627] <= r_data[27626];
                
                r_data[27628] <= r_data[27627];
                
                r_data[27629] <= r_data[27628];
                
                r_data[27630] <= r_data[27629];
                
                r_data[27631] <= r_data[27630];
                
                r_data[27632] <= r_data[27631];
                
                r_data[27633] <= r_data[27632];
                
                r_data[27634] <= r_data[27633];
                
                r_data[27635] <= r_data[27634];
                
                r_data[27636] <= r_data[27635];
                
                r_data[27637] <= r_data[27636];
                
                r_data[27638] <= r_data[27637];
                
                r_data[27639] <= r_data[27638];
                
                r_data[27640] <= r_data[27639];
                
                r_data[27641] <= r_data[27640];
                
                r_data[27642] <= r_data[27641];
                
                r_data[27643] <= r_data[27642];
                
                r_data[27644] <= r_data[27643];
                
                r_data[27645] <= r_data[27644];
                
                r_data[27646] <= r_data[27645];
                
                r_data[27647] <= r_data[27646];
                
                r_data[27648] <= r_data[27647];
                
                r_data[27649] <= r_data[27648];
                
                r_data[27650] <= r_data[27649];
                
                r_data[27651] <= r_data[27650];
                
                r_data[27652] <= r_data[27651];
                
                r_data[27653] <= r_data[27652];
                
                r_data[27654] <= r_data[27653];
                
                r_data[27655] <= r_data[27654];
                
                r_data[27656] <= r_data[27655];
                
                r_data[27657] <= r_data[27656];
                
                r_data[27658] <= r_data[27657];
                
                r_data[27659] <= r_data[27658];
                
                r_data[27660] <= r_data[27659];
                
                r_data[27661] <= r_data[27660];
                
                r_data[27662] <= r_data[27661];
                
                r_data[27663] <= r_data[27662];
                
                r_data[27664] <= r_data[27663];
                
                r_data[27665] <= r_data[27664];
                
                r_data[27666] <= r_data[27665];
                
                r_data[27667] <= r_data[27666];
                
                r_data[27668] <= r_data[27667];
                
                r_data[27669] <= r_data[27668];
                
                r_data[27670] <= r_data[27669];
                
                r_data[27671] <= r_data[27670];
                
                r_data[27672] <= r_data[27671];
                
                r_data[27673] <= r_data[27672];
                
                r_data[27674] <= r_data[27673];
                
                r_data[27675] <= r_data[27674];
                
                r_data[27676] <= r_data[27675];
                
                r_data[27677] <= r_data[27676];
                
                r_data[27678] <= r_data[27677];
                
                r_data[27679] <= r_data[27678];
                
                r_data[27680] <= r_data[27679];
                
                r_data[27681] <= r_data[27680];
                
                r_data[27682] <= r_data[27681];
                
                r_data[27683] <= r_data[27682];
                
                r_data[27684] <= r_data[27683];
                
                r_data[27685] <= r_data[27684];
                
                r_data[27686] <= r_data[27685];
                
                r_data[27687] <= r_data[27686];
                
                r_data[27688] <= r_data[27687];
                
                r_data[27689] <= r_data[27688];
                
                r_data[27690] <= r_data[27689];
                
                r_data[27691] <= r_data[27690];
                
                r_data[27692] <= r_data[27691];
                
                r_data[27693] <= r_data[27692];
                
                r_data[27694] <= r_data[27693];
                
                r_data[27695] <= r_data[27694];
                
                r_data[27696] <= r_data[27695];
                
                r_data[27697] <= r_data[27696];
                
                r_data[27698] <= r_data[27697];
                
                r_data[27699] <= r_data[27698];
                
                r_data[27700] <= r_data[27699];
                
                r_data[27701] <= r_data[27700];
                
                r_data[27702] <= r_data[27701];
                
                r_data[27703] <= r_data[27702];
                
                r_data[27704] <= r_data[27703];
                
                r_data[27705] <= r_data[27704];
                
                r_data[27706] <= r_data[27705];
                
                r_data[27707] <= r_data[27706];
                
                r_data[27708] <= r_data[27707];
                
                r_data[27709] <= r_data[27708];
                
                r_data[27710] <= r_data[27709];
                
                r_data[27711] <= r_data[27710];
                
                r_data[27712] <= r_data[27711];
                
                r_data[27713] <= r_data[27712];
                
                r_data[27714] <= r_data[27713];
                
                r_data[27715] <= r_data[27714];
                
                r_data[27716] <= r_data[27715];
                
                r_data[27717] <= r_data[27716];
                
                r_data[27718] <= r_data[27717];
                
                r_data[27719] <= r_data[27718];
                
                r_data[27720] <= r_data[27719];
                
                r_data[27721] <= r_data[27720];
                
                r_data[27722] <= r_data[27721];
                
                r_data[27723] <= r_data[27722];
                
                r_data[27724] <= r_data[27723];
                
                r_data[27725] <= r_data[27724];
                
                r_data[27726] <= r_data[27725];
                
                r_data[27727] <= r_data[27726];
                
                r_data[27728] <= r_data[27727];
                
                r_data[27729] <= r_data[27728];
                
                r_data[27730] <= r_data[27729];
                
                r_data[27731] <= r_data[27730];
                
                r_data[27732] <= r_data[27731];
                
                r_data[27733] <= r_data[27732];
                
                r_data[27734] <= r_data[27733];
                
                r_data[27735] <= r_data[27734];
                
                r_data[27736] <= r_data[27735];
                
                r_data[27737] <= r_data[27736];
                
                r_data[27738] <= r_data[27737];
                
                r_data[27739] <= r_data[27738];
                
                r_data[27740] <= r_data[27739];
                
                r_data[27741] <= r_data[27740];
                
                r_data[27742] <= r_data[27741];
                
                r_data[27743] <= r_data[27742];
                
                r_data[27744] <= r_data[27743];
                
                r_data[27745] <= r_data[27744];
                
                r_data[27746] <= r_data[27745];
                
                r_data[27747] <= r_data[27746];
                
                r_data[27748] <= r_data[27747];
                
                r_data[27749] <= r_data[27748];
                
                r_data[27750] <= r_data[27749];
                
                r_data[27751] <= r_data[27750];
                
                r_data[27752] <= r_data[27751];
                
                r_data[27753] <= r_data[27752];
                
                r_data[27754] <= r_data[27753];
                
                r_data[27755] <= r_data[27754];
                
                r_data[27756] <= r_data[27755];
                
                r_data[27757] <= r_data[27756];
                
                r_data[27758] <= r_data[27757];
                
                r_data[27759] <= r_data[27758];
                
                r_data[27760] <= r_data[27759];
                
                r_data[27761] <= r_data[27760];
                
                r_data[27762] <= r_data[27761];
                
                r_data[27763] <= r_data[27762];
                
                r_data[27764] <= r_data[27763];
                
                r_data[27765] <= r_data[27764];
                
                r_data[27766] <= r_data[27765];
                
                r_data[27767] <= r_data[27766];
                
                r_data[27768] <= r_data[27767];
                
                r_data[27769] <= r_data[27768];
                
                r_data[27770] <= r_data[27769];
                
                r_data[27771] <= r_data[27770];
                
                r_data[27772] <= r_data[27771];
                
                r_data[27773] <= r_data[27772];
                
                r_data[27774] <= r_data[27773];
                
                r_data[27775] <= r_data[27774];
                
                r_data[27776] <= r_data[27775];
                
                r_data[27777] <= r_data[27776];
                
                r_data[27778] <= r_data[27777];
                
                r_data[27779] <= r_data[27778];
                
                r_data[27780] <= r_data[27779];
                
                r_data[27781] <= r_data[27780];
                
                r_data[27782] <= r_data[27781];
                
                r_data[27783] <= r_data[27782];
                
                r_data[27784] <= r_data[27783];
                
                r_data[27785] <= r_data[27784];
                
                r_data[27786] <= r_data[27785];
                
                r_data[27787] <= r_data[27786];
                
                r_data[27788] <= r_data[27787];
                
                r_data[27789] <= r_data[27788];
                
                r_data[27790] <= r_data[27789];
                
                r_data[27791] <= r_data[27790];
                
                r_data[27792] <= r_data[27791];
                
                r_data[27793] <= r_data[27792];
                
                r_data[27794] <= r_data[27793];
                
                r_data[27795] <= r_data[27794];
                
                r_data[27796] <= r_data[27795];
                
                r_data[27797] <= r_data[27796];
                
                r_data[27798] <= r_data[27797];
                
                r_data[27799] <= r_data[27798];
                
                r_data[27800] <= r_data[27799];
                
                r_data[27801] <= r_data[27800];
                
                r_data[27802] <= r_data[27801];
                
                r_data[27803] <= r_data[27802];
                
                r_data[27804] <= r_data[27803];
                
                r_data[27805] <= r_data[27804];
                
                r_data[27806] <= r_data[27805];
                
                r_data[27807] <= r_data[27806];
                
                r_data[27808] <= r_data[27807];
                
                r_data[27809] <= r_data[27808];
                
                r_data[27810] <= r_data[27809];
                
                r_data[27811] <= r_data[27810];
                
                r_data[27812] <= r_data[27811];
                
                r_data[27813] <= r_data[27812];
                
                r_data[27814] <= r_data[27813];
                
                r_data[27815] <= r_data[27814];
                
                r_data[27816] <= r_data[27815];
                
                r_data[27817] <= r_data[27816];
                
                r_data[27818] <= r_data[27817];
                
                r_data[27819] <= r_data[27818];
                
                r_data[27820] <= r_data[27819];
                
                r_data[27821] <= r_data[27820];
                
                r_data[27822] <= r_data[27821];
                
                r_data[27823] <= r_data[27822];
                
                r_data[27824] <= r_data[27823];
                
                r_data[27825] <= r_data[27824];
                
                r_data[27826] <= r_data[27825];
                
                r_data[27827] <= r_data[27826];
                
                r_data[27828] <= r_data[27827];
                
                r_data[27829] <= r_data[27828];
                
                r_data[27830] <= r_data[27829];
                
                r_data[27831] <= r_data[27830];
                
                r_data[27832] <= r_data[27831];
                
                r_data[27833] <= r_data[27832];
                
                r_data[27834] <= r_data[27833];
                
                r_data[27835] <= r_data[27834];
                
                r_data[27836] <= r_data[27835];
                
                r_data[27837] <= r_data[27836];
                
                r_data[27838] <= r_data[27837];
                
                r_data[27839] <= r_data[27838];
                
                r_data[27840] <= r_data[27839];
                
                r_data[27841] <= r_data[27840];
                
                r_data[27842] <= r_data[27841];
                
                r_data[27843] <= r_data[27842];
                
                r_data[27844] <= r_data[27843];
                
                r_data[27845] <= r_data[27844];
                
                r_data[27846] <= r_data[27845];
                
                r_data[27847] <= r_data[27846];
                
                r_data[27848] <= r_data[27847];
                
                r_data[27849] <= r_data[27848];
                
                r_data[27850] <= r_data[27849];
                
                r_data[27851] <= r_data[27850];
                
                r_data[27852] <= r_data[27851];
                
                r_data[27853] <= r_data[27852];
                
                r_data[27854] <= r_data[27853];
                
                r_data[27855] <= r_data[27854];
                
                r_data[27856] <= r_data[27855];
                
                r_data[27857] <= r_data[27856];
                
                r_data[27858] <= r_data[27857];
                
                r_data[27859] <= r_data[27858];
                
                r_data[27860] <= r_data[27859];
                
                r_data[27861] <= r_data[27860];
                
                r_data[27862] <= r_data[27861];
                
                r_data[27863] <= r_data[27862];
                
                r_data[27864] <= r_data[27863];
                
                r_data[27865] <= r_data[27864];
                
                r_data[27866] <= r_data[27865];
                
                r_data[27867] <= r_data[27866];
                
                r_data[27868] <= r_data[27867];
                
                r_data[27869] <= r_data[27868];
                
                r_data[27870] <= r_data[27869];
                
                r_data[27871] <= r_data[27870];
                
                r_data[27872] <= r_data[27871];
                
                r_data[27873] <= r_data[27872];
                
                r_data[27874] <= r_data[27873];
                
                r_data[27875] <= r_data[27874];
                
                r_data[27876] <= r_data[27875];
                
                r_data[27877] <= r_data[27876];
                
                r_data[27878] <= r_data[27877];
                
                r_data[27879] <= r_data[27878];
                
                r_data[27880] <= r_data[27879];
                
                r_data[27881] <= r_data[27880];
                
                r_data[27882] <= r_data[27881];
                
                r_data[27883] <= r_data[27882];
                
                r_data[27884] <= r_data[27883];
                
                r_data[27885] <= r_data[27884];
                
                r_data[27886] <= r_data[27885];
                
                r_data[27887] <= r_data[27886];
                
                r_data[27888] <= r_data[27887];
                
                r_data[27889] <= r_data[27888];
                
                r_data[27890] <= r_data[27889];
                
                r_data[27891] <= r_data[27890];
                
                r_data[27892] <= r_data[27891];
                
                r_data[27893] <= r_data[27892];
                
                r_data[27894] <= r_data[27893];
                
                r_data[27895] <= r_data[27894];
                
                r_data[27896] <= r_data[27895];
                
                r_data[27897] <= r_data[27896];
                
                r_data[27898] <= r_data[27897];
                
                r_data[27899] <= r_data[27898];
                
                r_data[27900] <= r_data[27899];
                
                r_data[27901] <= r_data[27900];
                
                r_data[27902] <= r_data[27901];
                
                r_data[27903] <= r_data[27902];
                
                r_data[27904] <= r_data[27903];
                
                r_data[27905] <= r_data[27904];
                
                r_data[27906] <= r_data[27905];
                
                r_data[27907] <= r_data[27906];
                
                r_data[27908] <= r_data[27907];
                
                r_data[27909] <= r_data[27908];
                
                r_data[27910] <= r_data[27909];
                
                r_data[27911] <= r_data[27910];
                
                r_data[27912] <= r_data[27911];
                
                r_data[27913] <= r_data[27912];
                
                r_data[27914] <= r_data[27913];
                
                r_data[27915] <= r_data[27914];
                
                r_data[27916] <= r_data[27915];
                
                r_data[27917] <= r_data[27916];
                
                r_data[27918] <= r_data[27917];
                
                r_data[27919] <= r_data[27918];
                
                r_data[27920] <= r_data[27919];
                
                r_data[27921] <= r_data[27920];
                
                r_data[27922] <= r_data[27921];
                
                r_data[27923] <= r_data[27922];
                
                r_data[27924] <= r_data[27923];
                
                r_data[27925] <= r_data[27924];
                
                r_data[27926] <= r_data[27925];
                
                r_data[27927] <= r_data[27926];
                
                r_data[27928] <= r_data[27927];
                
                r_data[27929] <= r_data[27928];
                
                r_data[27930] <= r_data[27929];
                
                r_data[27931] <= r_data[27930];
                
                r_data[27932] <= r_data[27931];
                
                r_data[27933] <= r_data[27932];
                
                r_data[27934] <= r_data[27933];
                
                r_data[27935] <= r_data[27934];
                
                r_data[27936] <= r_data[27935];
                
                r_data[27937] <= r_data[27936];
                
                r_data[27938] <= r_data[27937];
                
                r_data[27939] <= r_data[27938];
                
                r_data[27940] <= r_data[27939];
                
                r_data[27941] <= r_data[27940];
                
                r_data[27942] <= r_data[27941];
                
                r_data[27943] <= r_data[27942];
                
                r_data[27944] <= r_data[27943];
                
                r_data[27945] <= r_data[27944];
                
                r_data[27946] <= r_data[27945];
                
                r_data[27947] <= r_data[27946];
                
                r_data[27948] <= r_data[27947];
                
                r_data[27949] <= r_data[27948];
                
                r_data[27950] <= r_data[27949];
                
                r_data[27951] <= r_data[27950];
                
                r_data[27952] <= r_data[27951];
                
                r_data[27953] <= r_data[27952];
                
                r_data[27954] <= r_data[27953];
                
                r_data[27955] <= r_data[27954];
                
                r_data[27956] <= r_data[27955];
                
                r_data[27957] <= r_data[27956];
                
                r_data[27958] <= r_data[27957];
                
                r_data[27959] <= r_data[27958];
                
                r_data[27960] <= r_data[27959];
                
                r_data[27961] <= r_data[27960];
                
                r_data[27962] <= r_data[27961];
                
                r_data[27963] <= r_data[27962];
                
                r_data[27964] <= r_data[27963];
                
                r_data[27965] <= r_data[27964];
                
                r_data[27966] <= r_data[27965];
                
                r_data[27967] <= r_data[27966];
                
                r_data[27968] <= r_data[27967];
                
                r_data[27969] <= r_data[27968];
                
                r_data[27970] <= r_data[27969];
                
                r_data[27971] <= r_data[27970];
                
                r_data[27972] <= r_data[27971];
                
                r_data[27973] <= r_data[27972];
                
                r_data[27974] <= r_data[27973];
                
                r_data[27975] <= r_data[27974];
                
                r_data[27976] <= r_data[27975];
                
                r_data[27977] <= r_data[27976];
                
                r_data[27978] <= r_data[27977];
                
                r_data[27979] <= r_data[27978];
                
                r_data[27980] <= r_data[27979];
                
                r_data[27981] <= r_data[27980];
                
                r_data[27982] <= r_data[27981];
                
                r_data[27983] <= r_data[27982];
                
                r_data[27984] <= r_data[27983];
                
                r_data[27985] <= r_data[27984];
                
                r_data[27986] <= r_data[27985];
                
                r_data[27987] <= r_data[27986];
                
                r_data[27988] <= r_data[27987];
                
                r_data[27989] <= r_data[27988];
                
                r_data[27990] <= r_data[27989];
                
                r_data[27991] <= r_data[27990];
                
                r_data[27992] <= r_data[27991];
                
                r_data[27993] <= r_data[27992];
                
                r_data[27994] <= r_data[27993];
                
                r_data[27995] <= r_data[27994];
                
                r_data[27996] <= r_data[27995];
                
                r_data[27997] <= r_data[27996];
                
                r_data[27998] <= r_data[27997];
                
                r_data[27999] <= r_data[27998];
                
                r_data[28000] <= r_data[27999];
                
                r_data[28001] <= r_data[28000];
                
                r_data[28002] <= r_data[28001];
                
                r_data[28003] <= r_data[28002];
                
                r_data[28004] <= r_data[28003];
                
                r_data[28005] <= r_data[28004];
                
                r_data[28006] <= r_data[28005];
                
                r_data[28007] <= r_data[28006];
                
                r_data[28008] <= r_data[28007];
                
                r_data[28009] <= r_data[28008];
                
                r_data[28010] <= r_data[28009];
                
                r_data[28011] <= r_data[28010];
                
                r_data[28012] <= r_data[28011];
                
                r_data[28013] <= r_data[28012];
                
                r_data[28014] <= r_data[28013];
                
                r_data[28015] <= r_data[28014];
                
                r_data[28016] <= r_data[28015];
                
                r_data[28017] <= r_data[28016];
                
                r_data[28018] <= r_data[28017];
                
                r_data[28019] <= r_data[28018];
                
                r_data[28020] <= r_data[28019];
                
                r_data[28021] <= r_data[28020];
                
                r_data[28022] <= r_data[28021];
                
                r_data[28023] <= r_data[28022];
                
                r_data[28024] <= r_data[28023];
                
                r_data[28025] <= r_data[28024];
                
                r_data[28026] <= r_data[28025];
                
                r_data[28027] <= r_data[28026];
                
                r_data[28028] <= r_data[28027];
                
                r_data[28029] <= r_data[28028];
                
                r_data[28030] <= r_data[28029];
                
                r_data[28031] <= r_data[28030];
                
                r_data[28032] <= r_data[28031];
                
                r_data[28033] <= r_data[28032];
                
                r_data[28034] <= r_data[28033];
                
                r_data[28035] <= r_data[28034];
                
                r_data[28036] <= r_data[28035];
                
                r_data[28037] <= r_data[28036];
                
                r_data[28038] <= r_data[28037];
                
                r_data[28039] <= r_data[28038];
                
                r_data[28040] <= r_data[28039];
                
                r_data[28041] <= r_data[28040];
                
                r_data[28042] <= r_data[28041];
                
                r_data[28043] <= r_data[28042];
                
                r_data[28044] <= r_data[28043];
                
                r_data[28045] <= r_data[28044];
                
                r_data[28046] <= r_data[28045];
                
                r_data[28047] <= r_data[28046];
                
                r_data[28048] <= r_data[28047];
                
                r_data[28049] <= r_data[28048];
                
                r_data[28050] <= r_data[28049];
                
                r_data[28051] <= r_data[28050];
                
                r_data[28052] <= r_data[28051];
                
                r_data[28053] <= r_data[28052];
                
                r_data[28054] <= r_data[28053];
                
                r_data[28055] <= r_data[28054];
                
                r_data[28056] <= r_data[28055];
                
                r_data[28057] <= r_data[28056];
                
                r_data[28058] <= r_data[28057];
                
                r_data[28059] <= r_data[28058];
                
                r_data[28060] <= r_data[28059];
                
                r_data[28061] <= r_data[28060];
                
                r_data[28062] <= r_data[28061];
                
                r_data[28063] <= r_data[28062];
                
                r_data[28064] <= r_data[28063];
                
                r_data[28065] <= r_data[28064];
                
                r_data[28066] <= r_data[28065];
                
                r_data[28067] <= r_data[28066];
                
                r_data[28068] <= r_data[28067];
                
                r_data[28069] <= r_data[28068];
                
                r_data[28070] <= r_data[28069];
                
                r_data[28071] <= r_data[28070];
                
                r_data[28072] <= r_data[28071];
                
                r_data[28073] <= r_data[28072];
                
                r_data[28074] <= r_data[28073];
                
                r_data[28075] <= r_data[28074];
                
                r_data[28076] <= r_data[28075];
                
                r_data[28077] <= r_data[28076];
                
                r_data[28078] <= r_data[28077];
                
                r_data[28079] <= r_data[28078];
                
                r_data[28080] <= r_data[28079];
                
                r_data[28081] <= r_data[28080];
                
                r_data[28082] <= r_data[28081];
                
                r_data[28083] <= r_data[28082];
                
                r_data[28084] <= r_data[28083];
                
                r_data[28085] <= r_data[28084];
                
                r_data[28086] <= r_data[28085];
                
                r_data[28087] <= r_data[28086];
                
                r_data[28088] <= r_data[28087];
                
                r_data[28089] <= r_data[28088];
                
                r_data[28090] <= r_data[28089];
                
                r_data[28091] <= r_data[28090];
                
                r_data[28092] <= r_data[28091];
                
                r_data[28093] <= r_data[28092];
                
                r_data[28094] <= r_data[28093];
                
                r_data[28095] <= r_data[28094];
                
                r_data[28096] <= r_data[28095];
                
                r_data[28097] <= r_data[28096];
                
                r_data[28098] <= r_data[28097];
                
                r_data[28099] <= r_data[28098];
                
                r_data[28100] <= r_data[28099];
                
                r_data[28101] <= r_data[28100];
                
                r_data[28102] <= r_data[28101];
                
                r_data[28103] <= r_data[28102];
                
                r_data[28104] <= r_data[28103];
                
                r_data[28105] <= r_data[28104];
                
                r_data[28106] <= r_data[28105];
                
                r_data[28107] <= r_data[28106];
                
                r_data[28108] <= r_data[28107];
                
                r_data[28109] <= r_data[28108];
                
                r_data[28110] <= r_data[28109];
                
                r_data[28111] <= r_data[28110];
                
                r_data[28112] <= r_data[28111];
                
                r_data[28113] <= r_data[28112];
                
                r_data[28114] <= r_data[28113];
                
                r_data[28115] <= r_data[28114];
                
                r_data[28116] <= r_data[28115];
                
                r_data[28117] <= r_data[28116];
                
                r_data[28118] <= r_data[28117];
                
                r_data[28119] <= r_data[28118];
                
                r_data[28120] <= r_data[28119];
                
                r_data[28121] <= r_data[28120];
                
                r_data[28122] <= r_data[28121];
                
                r_data[28123] <= r_data[28122];
                
                r_data[28124] <= r_data[28123];
                
                r_data[28125] <= r_data[28124];
                
                r_data[28126] <= r_data[28125];
                
                r_data[28127] <= r_data[28126];
                
                r_data[28128] <= r_data[28127];
                
                r_data[28129] <= r_data[28128];
                
                r_data[28130] <= r_data[28129];
                
                r_data[28131] <= r_data[28130];
                
                r_data[28132] <= r_data[28131];
                
                r_data[28133] <= r_data[28132];
                
                r_data[28134] <= r_data[28133];
                
                r_data[28135] <= r_data[28134];
                
                r_data[28136] <= r_data[28135];
                
                r_data[28137] <= r_data[28136];
                
                r_data[28138] <= r_data[28137];
                
                r_data[28139] <= r_data[28138];
                
                r_data[28140] <= r_data[28139];
                
                r_data[28141] <= r_data[28140];
                
                r_data[28142] <= r_data[28141];
                
                r_data[28143] <= r_data[28142];
                
                r_data[28144] <= r_data[28143];
                
                r_data[28145] <= r_data[28144];
                
                r_data[28146] <= r_data[28145];
                
                r_data[28147] <= r_data[28146];
                
                r_data[28148] <= r_data[28147];
                
                r_data[28149] <= r_data[28148];
                
                r_data[28150] <= r_data[28149];
                
                r_data[28151] <= r_data[28150];
                
                r_data[28152] <= r_data[28151];
                
                r_data[28153] <= r_data[28152];
                
                r_data[28154] <= r_data[28153];
                
                r_data[28155] <= r_data[28154];
                
                r_data[28156] <= r_data[28155];
                
                r_data[28157] <= r_data[28156];
                
                r_data[28158] <= r_data[28157];
                
                r_data[28159] <= r_data[28158];
                
                r_data[28160] <= r_data[28159];
                
                r_data[28161] <= r_data[28160];
                
                r_data[28162] <= r_data[28161];
                
                r_data[28163] <= r_data[28162];
                
                r_data[28164] <= r_data[28163];
                
                r_data[28165] <= r_data[28164];
                
                r_data[28166] <= r_data[28165];
                
                r_data[28167] <= r_data[28166];
                
                r_data[28168] <= r_data[28167];
                
                r_data[28169] <= r_data[28168];
                
                r_data[28170] <= r_data[28169];
                
                r_data[28171] <= r_data[28170];
                
                r_data[28172] <= r_data[28171];
                
                r_data[28173] <= r_data[28172];
                
                r_data[28174] <= r_data[28173];
                
                r_data[28175] <= r_data[28174];
                
                r_data[28176] <= r_data[28175];
                
                r_data[28177] <= r_data[28176];
                
                r_data[28178] <= r_data[28177];
                
                r_data[28179] <= r_data[28178];
                
                r_data[28180] <= r_data[28179];
                
                r_data[28181] <= r_data[28180];
                
                r_data[28182] <= r_data[28181];
                
                r_data[28183] <= r_data[28182];
                
                r_data[28184] <= r_data[28183];
                
                r_data[28185] <= r_data[28184];
                
                r_data[28186] <= r_data[28185];
                
                r_data[28187] <= r_data[28186];
                
                r_data[28188] <= r_data[28187];
                
                r_data[28189] <= r_data[28188];
                
                r_data[28190] <= r_data[28189];
                
                r_data[28191] <= r_data[28190];
                
                r_data[28192] <= r_data[28191];
                
                r_data[28193] <= r_data[28192];
                
                r_data[28194] <= r_data[28193];
                
                r_data[28195] <= r_data[28194];
                
                r_data[28196] <= r_data[28195];
                
                r_data[28197] <= r_data[28196];
                
                r_data[28198] <= r_data[28197];
                
                r_data[28199] <= r_data[28198];
                
                r_data[28200] <= r_data[28199];
                
                r_data[28201] <= r_data[28200];
                
                r_data[28202] <= r_data[28201];
                
                r_data[28203] <= r_data[28202];
                
                r_data[28204] <= r_data[28203];
                
                r_data[28205] <= r_data[28204];
                
                r_data[28206] <= r_data[28205];
                
                r_data[28207] <= r_data[28206];
                
                r_data[28208] <= r_data[28207];
                
                r_data[28209] <= r_data[28208];
                
                r_data[28210] <= r_data[28209];
                
                r_data[28211] <= r_data[28210];
                
                r_data[28212] <= r_data[28211];
                
                r_data[28213] <= r_data[28212];
                
                r_data[28214] <= r_data[28213];
                
                r_data[28215] <= r_data[28214];
                
                r_data[28216] <= r_data[28215];
                
                r_data[28217] <= r_data[28216];
                
                r_data[28218] <= r_data[28217];
                
                r_data[28219] <= r_data[28218];
                
                r_data[28220] <= r_data[28219];
                
                r_data[28221] <= r_data[28220];
                
                r_data[28222] <= r_data[28221];
                
                r_data[28223] <= r_data[28222];
                
                r_data[28224] <= r_data[28223];
                
                r_data[28225] <= r_data[28224];
                
                r_data[28226] <= r_data[28225];
                
                r_data[28227] <= r_data[28226];
                
                r_data[28228] <= r_data[28227];
                
                r_data[28229] <= r_data[28228];
                
                r_data[28230] <= r_data[28229];
                
                r_data[28231] <= r_data[28230];
                
                r_data[28232] <= r_data[28231];
                
                r_data[28233] <= r_data[28232];
                
                r_data[28234] <= r_data[28233];
                
                r_data[28235] <= r_data[28234];
                
                r_data[28236] <= r_data[28235];
                
                r_data[28237] <= r_data[28236];
                
                r_data[28238] <= r_data[28237];
                
                r_data[28239] <= r_data[28238];
                
                r_data[28240] <= r_data[28239];
                
                r_data[28241] <= r_data[28240];
                
                r_data[28242] <= r_data[28241];
                
                r_data[28243] <= r_data[28242];
                
                r_data[28244] <= r_data[28243];
                
                r_data[28245] <= r_data[28244];
                
                r_data[28246] <= r_data[28245];
                
                r_data[28247] <= r_data[28246];
                
                r_data[28248] <= r_data[28247];
                
                r_data[28249] <= r_data[28248];
                
                r_data[28250] <= r_data[28249];
                
                r_data[28251] <= r_data[28250];
                
                r_data[28252] <= r_data[28251];
                
                r_data[28253] <= r_data[28252];
                
                r_data[28254] <= r_data[28253];
                
                r_data[28255] <= r_data[28254];
                
                r_data[28256] <= r_data[28255];
                
                r_data[28257] <= r_data[28256];
                
                r_data[28258] <= r_data[28257];
                
                r_data[28259] <= r_data[28258];
                
                r_data[28260] <= r_data[28259];
                
                r_data[28261] <= r_data[28260];
                
                r_data[28262] <= r_data[28261];
                
                r_data[28263] <= r_data[28262];
                
                r_data[28264] <= r_data[28263];
                
                r_data[28265] <= r_data[28264];
                
                r_data[28266] <= r_data[28265];
                
                r_data[28267] <= r_data[28266];
                
                r_data[28268] <= r_data[28267];
                
                r_data[28269] <= r_data[28268];
                
                r_data[28270] <= r_data[28269];
                
                r_data[28271] <= r_data[28270];
                
                r_data[28272] <= r_data[28271];
                
                r_data[28273] <= r_data[28272];
                
                r_data[28274] <= r_data[28273];
                
                r_data[28275] <= r_data[28274];
                
                r_data[28276] <= r_data[28275];
                
                r_data[28277] <= r_data[28276];
                
                r_data[28278] <= r_data[28277];
                
                r_data[28279] <= r_data[28278];
                
                r_data[28280] <= r_data[28279];
                
                r_data[28281] <= r_data[28280];
                
                r_data[28282] <= r_data[28281];
                
                r_data[28283] <= r_data[28282];
                
                r_data[28284] <= r_data[28283];
                
                r_data[28285] <= r_data[28284];
                
                r_data[28286] <= r_data[28285];
                
                r_data[28287] <= r_data[28286];
                
                r_data[28288] <= r_data[28287];
                
                r_data[28289] <= r_data[28288];
                
                r_data[28290] <= r_data[28289];
                
                r_data[28291] <= r_data[28290];
                
                r_data[28292] <= r_data[28291];
                
                r_data[28293] <= r_data[28292];
                
                r_data[28294] <= r_data[28293];
                
                r_data[28295] <= r_data[28294];
                
                r_data[28296] <= r_data[28295];
                
                r_data[28297] <= r_data[28296];
                
                r_data[28298] <= r_data[28297];
                
                r_data[28299] <= r_data[28298];
                
                r_data[28300] <= r_data[28299];
                
                r_data[28301] <= r_data[28300];
                
                r_data[28302] <= r_data[28301];
                
                r_data[28303] <= r_data[28302];
                
                r_data[28304] <= r_data[28303];
                
                r_data[28305] <= r_data[28304];
                
                r_data[28306] <= r_data[28305];
                
                r_data[28307] <= r_data[28306];
                
                r_data[28308] <= r_data[28307];
                
                r_data[28309] <= r_data[28308];
                
                r_data[28310] <= r_data[28309];
                
                r_data[28311] <= r_data[28310];
                
                r_data[28312] <= r_data[28311];
                
                r_data[28313] <= r_data[28312];
                
                r_data[28314] <= r_data[28313];
                
                r_data[28315] <= r_data[28314];
                
                r_data[28316] <= r_data[28315];
                
                r_data[28317] <= r_data[28316];
                
                r_data[28318] <= r_data[28317];
                
                r_data[28319] <= r_data[28318];
                
                r_data[28320] <= r_data[28319];
                
                r_data[28321] <= r_data[28320];
                
                r_data[28322] <= r_data[28321];
                
                r_data[28323] <= r_data[28322];
                
                r_data[28324] <= r_data[28323];
                
                r_data[28325] <= r_data[28324];
                
                r_data[28326] <= r_data[28325];
                
                r_data[28327] <= r_data[28326];
                
                r_data[28328] <= r_data[28327];
                
                r_data[28329] <= r_data[28328];
                
                r_data[28330] <= r_data[28329];
                
                r_data[28331] <= r_data[28330];
                
                r_data[28332] <= r_data[28331];
                
                r_data[28333] <= r_data[28332];
                
                r_data[28334] <= r_data[28333];
                
                r_data[28335] <= r_data[28334];
                
                r_data[28336] <= r_data[28335];
                
                r_data[28337] <= r_data[28336];
                
                r_data[28338] <= r_data[28337];
                
                r_data[28339] <= r_data[28338];
                
                r_data[28340] <= r_data[28339];
                
                r_data[28341] <= r_data[28340];
                
                r_data[28342] <= r_data[28341];
                
                r_data[28343] <= r_data[28342];
                
                r_data[28344] <= r_data[28343];
                
                r_data[28345] <= r_data[28344];
                
                r_data[28346] <= r_data[28345];
                
                r_data[28347] <= r_data[28346];
                
                r_data[28348] <= r_data[28347];
                
                r_data[28349] <= r_data[28348];
                
                r_data[28350] <= r_data[28349];
                
                r_data[28351] <= r_data[28350];
                
                r_data[28352] <= r_data[28351];
                
                r_data[28353] <= r_data[28352];
                
                r_data[28354] <= r_data[28353];
                
                r_data[28355] <= r_data[28354];
                
                r_data[28356] <= r_data[28355];
                
                r_data[28357] <= r_data[28356];
                
                r_data[28358] <= r_data[28357];
                
                r_data[28359] <= r_data[28358];
                
                r_data[28360] <= r_data[28359];
                
                r_data[28361] <= r_data[28360];
                
                r_data[28362] <= r_data[28361];
                
                r_data[28363] <= r_data[28362];
                
                r_data[28364] <= r_data[28363];
                
                r_data[28365] <= r_data[28364];
                
                r_data[28366] <= r_data[28365];
                
                r_data[28367] <= r_data[28366];
                
                r_data[28368] <= r_data[28367];
                
                r_data[28369] <= r_data[28368];
                
                r_data[28370] <= r_data[28369];
                
                r_data[28371] <= r_data[28370];
                
                r_data[28372] <= r_data[28371];
                
                r_data[28373] <= r_data[28372];
                
                r_data[28374] <= r_data[28373];
                
                r_data[28375] <= r_data[28374];
                
                r_data[28376] <= r_data[28375];
                
                r_data[28377] <= r_data[28376];
                
                r_data[28378] <= r_data[28377];
                
                r_data[28379] <= r_data[28378];
                
                r_data[28380] <= r_data[28379];
                
                r_data[28381] <= r_data[28380];
                
                r_data[28382] <= r_data[28381];
                
                r_data[28383] <= r_data[28382];
                
                r_data[28384] <= r_data[28383];
                
                r_data[28385] <= r_data[28384];
                
                r_data[28386] <= r_data[28385];
                
                r_data[28387] <= r_data[28386];
                
                r_data[28388] <= r_data[28387];
                
                r_data[28389] <= r_data[28388];
                
                r_data[28390] <= r_data[28389];
                
                r_data[28391] <= r_data[28390];
                
                r_data[28392] <= r_data[28391];
                
                r_data[28393] <= r_data[28392];
                
                r_data[28394] <= r_data[28393];
                
                r_data[28395] <= r_data[28394];
                
                r_data[28396] <= r_data[28395];
                
                r_data[28397] <= r_data[28396];
                
                r_data[28398] <= r_data[28397];
                
                r_data[28399] <= r_data[28398];
                
                r_data[28400] <= r_data[28399];
                
                r_data[28401] <= r_data[28400];
                
                r_data[28402] <= r_data[28401];
                
                r_data[28403] <= r_data[28402];
                
                r_data[28404] <= r_data[28403];
                
                r_data[28405] <= r_data[28404];
                
                r_data[28406] <= r_data[28405];
                
                r_data[28407] <= r_data[28406];
                
                r_data[28408] <= r_data[28407];
                
                r_data[28409] <= r_data[28408];
                
                r_data[28410] <= r_data[28409];
                
                r_data[28411] <= r_data[28410];
                
                r_data[28412] <= r_data[28411];
                
                r_data[28413] <= r_data[28412];
                
                r_data[28414] <= r_data[28413];
                
                r_data[28415] <= r_data[28414];
                
                r_data[28416] <= r_data[28415];
                
                r_data[28417] <= r_data[28416];
                
                r_data[28418] <= r_data[28417];
                
                r_data[28419] <= r_data[28418];
                
                r_data[28420] <= r_data[28419];
                
                r_data[28421] <= r_data[28420];
                
                r_data[28422] <= r_data[28421];
                
                r_data[28423] <= r_data[28422];
                
                r_data[28424] <= r_data[28423];
                
                r_data[28425] <= r_data[28424];
                
                r_data[28426] <= r_data[28425];
                
                r_data[28427] <= r_data[28426];
                
                r_data[28428] <= r_data[28427];
                
                r_data[28429] <= r_data[28428];
                
                r_data[28430] <= r_data[28429];
                
                r_data[28431] <= r_data[28430];
                
                r_data[28432] <= r_data[28431];
                
                r_data[28433] <= r_data[28432];
                
                r_data[28434] <= r_data[28433];
                
                r_data[28435] <= r_data[28434];
                
                r_data[28436] <= r_data[28435];
                
                r_data[28437] <= r_data[28436];
                
                r_data[28438] <= r_data[28437];
                
                r_data[28439] <= r_data[28438];
                
                r_data[28440] <= r_data[28439];
                
                r_data[28441] <= r_data[28440];
                
                r_data[28442] <= r_data[28441];
                
                r_data[28443] <= r_data[28442];
                
                r_data[28444] <= r_data[28443];
                
                r_data[28445] <= r_data[28444];
                
                r_data[28446] <= r_data[28445];
                
                r_data[28447] <= r_data[28446];
                
                r_data[28448] <= r_data[28447];
                
                r_data[28449] <= r_data[28448];
                
                r_data[28450] <= r_data[28449];
                
                r_data[28451] <= r_data[28450];
                
                r_data[28452] <= r_data[28451];
                
                r_data[28453] <= r_data[28452];
                
                r_data[28454] <= r_data[28453];
                
                r_data[28455] <= r_data[28454];
                
                r_data[28456] <= r_data[28455];
                
                r_data[28457] <= r_data[28456];
                
                r_data[28458] <= r_data[28457];
                
                r_data[28459] <= r_data[28458];
                
                r_data[28460] <= r_data[28459];
                
                r_data[28461] <= r_data[28460];
                
                r_data[28462] <= r_data[28461];
                
                r_data[28463] <= r_data[28462];
                
                r_data[28464] <= r_data[28463];
                
                r_data[28465] <= r_data[28464];
                
                r_data[28466] <= r_data[28465];
                
                r_data[28467] <= r_data[28466];
                
                r_data[28468] <= r_data[28467];
                
                r_data[28469] <= r_data[28468];
                
                r_data[28470] <= r_data[28469];
                
                r_data[28471] <= r_data[28470];
                
                r_data[28472] <= r_data[28471];
                
                r_data[28473] <= r_data[28472];
                
                r_data[28474] <= r_data[28473];
                
                r_data[28475] <= r_data[28474];
                
                r_data[28476] <= r_data[28475];
                
                r_data[28477] <= r_data[28476];
                
                r_data[28478] <= r_data[28477];
                
                r_data[28479] <= r_data[28478];
                
                r_data[28480] <= r_data[28479];
                
                r_data[28481] <= r_data[28480];
                
                r_data[28482] <= r_data[28481];
                
                r_data[28483] <= r_data[28482];
                
                r_data[28484] <= r_data[28483];
                
                r_data[28485] <= r_data[28484];
                
                r_data[28486] <= r_data[28485];
                
                r_data[28487] <= r_data[28486];
                
                r_data[28488] <= r_data[28487];
                
                r_data[28489] <= r_data[28488];
                
                r_data[28490] <= r_data[28489];
                
                r_data[28491] <= r_data[28490];
                
                r_data[28492] <= r_data[28491];
                
                r_data[28493] <= r_data[28492];
                
                r_data[28494] <= r_data[28493];
                
                r_data[28495] <= r_data[28494];
                
                r_data[28496] <= r_data[28495];
                
                r_data[28497] <= r_data[28496];
                
                r_data[28498] <= r_data[28497];
                
                r_data[28499] <= r_data[28498];
                
                r_data[28500] <= r_data[28499];
                
                r_data[28501] <= r_data[28500];
                
                r_data[28502] <= r_data[28501];
                
                r_data[28503] <= r_data[28502];
                
                r_data[28504] <= r_data[28503];
                
                r_data[28505] <= r_data[28504];
                
                r_data[28506] <= r_data[28505];
                
                r_data[28507] <= r_data[28506];
                
                r_data[28508] <= r_data[28507];
                
                r_data[28509] <= r_data[28508];
                
                r_data[28510] <= r_data[28509];
                
                r_data[28511] <= r_data[28510];
                
                r_data[28512] <= r_data[28511];
                
                r_data[28513] <= r_data[28512];
                
                r_data[28514] <= r_data[28513];
                
                r_data[28515] <= r_data[28514];
                
                r_data[28516] <= r_data[28515];
                
                r_data[28517] <= r_data[28516];
                
                r_data[28518] <= r_data[28517];
                
                r_data[28519] <= r_data[28518];
                
                r_data[28520] <= r_data[28519];
                
                r_data[28521] <= r_data[28520];
                
                r_data[28522] <= r_data[28521];
                
                r_data[28523] <= r_data[28522];
                
                r_data[28524] <= r_data[28523];
                
                r_data[28525] <= r_data[28524];
                
                r_data[28526] <= r_data[28525];
                
                r_data[28527] <= r_data[28526];
                
                r_data[28528] <= r_data[28527];
                
                r_data[28529] <= r_data[28528];
                
                r_data[28530] <= r_data[28529];
                
                r_data[28531] <= r_data[28530];
                
                r_data[28532] <= r_data[28531];
                
                r_data[28533] <= r_data[28532];
                
                r_data[28534] <= r_data[28533];
                
                r_data[28535] <= r_data[28534];
                
                r_data[28536] <= r_data[28535];
                
                r_data[28537] <= r_data[28536];
                
                r_data[28538] <= r_data[28537];
                
                r_data[28539] <= r_data[28538];
                
                r_data[28540] <= r_data[28539];
                
                r_data[28541] <= r_data[28540];
                
                r_data[28542] <= r_data[28541];
                
                r_data[28543] <= r_data[28542];
                
                r_data[28544] <= r_data[28543];
                
                r_data[28545] <= r_data[28544];
                
                r_data[28546] <= r_data[28545];
                
                r_data[28547] <= r_data[28546];
                
                r_data[28548] <= r_data[28547];
                
                r_data[28549] <= r_data[28548];
                
                r_data[28550] <= r_data[28549];
                
                r_data[28551] <= r_data[28550];
                
                r_data[28552] <= r_data[28551];
                
                r_data[28553] <= r_data[28552];
                
                r_data[28554] <= r_data[28553];
                
                r_data[28555] <= r_data[28554];
                
                r_data[28556] <= r_data[28555];
                
                r_data[28557] <= r_data[28556];
                
                r_data[28558] <= r_data[28557];
                
                r_data[28559] <= r_data[28558];
                
                r_data[28560] <= r_data[28559];
                
                r_data[28561] <= r_data[28560];
                
                r_data[28562] <= r_data[28561];
                
                r_data[28563] <= r_data[28562];
                
                r_data[28564] <= r_data[28563];
                
                r_data[28565] <= r_data[28564];
                
                r_data[28566] <= r_data[28565];
                
                r_data[28567] <= r_data[28566];
                
                r_data[28568] <= r_data[28567];
                
                r_data[28569] <= r_data[28568];
                
                r_data[28570] <= r_data[28569];
                
                r_data[28571] <= r_data[28570];
                
                r_data[28572] <= r_data[28571];
                
                r_data[28573] <= r_data[28572];
                
                r_data[28574] <= r_data[28573];
                
                r_data[28575] <= r_data[28574];
                
                r_data[28576] <= r_data[28575];
                
                r_data[28577] <= r_data[28576];
                
                r_data[28578] <= r_data[28577];
                
                r_data[28579] <= r_data[28578];
                
                r_data[28580] <= r_data[28579];
                
                r_data[28581] <= r_data[28580];
                
                r_data[28582] <= r_data[28581];
                
                r_data[28583] <= r_data[28582];
                
                r_data[28584] <= r_data[28583];
                
                r_data[28585] <= r_data[28584];
                
                r_data[28586] <= r_data[28585];
                
                r_data[28587] <= r_data[28586];
                
                r_data[28588] <= r_data[28587];
                
                r_data[28589] <= r_data[28588];
                
                r_data[28590] <= r_data[28589];
                
                r_data[28591] <= r_data[28590];
                
                r_data[28592] <= r_data[28591];
                
                r_data[28593] <= r_data[28592];
                
                r_data[28594] <= r_data[28593];
                
                r_data[28595] <= r_data[28594];
                
                r_data[28596] <= r_data[28595];
                
                r_data[28597] <= r_data[28596];
                
                r_data[28598] <= r_data[28597];
                
                r_data[28599] <= r_data[28598];
                
                r_data[28600] <= r_data[28599];
                
                r_data[28601] <= r_data[28600];
                
                r_data[28602] <= r_data[28601];
                
                r_data[28603] <= r_data[28602];
                
                r_data[28604] <= r_data[28603];
                
                r_data[28605] <= r_data[28604];
                
                r_data[28606] <= r_data[28605];
                
                r_data[28607] <= r_data[28606];
                
                r_data[28608] <= r_data[28607];
                
                r_data[28609] <= r_data[28608];
                
                r_data[28610] <= r_data[28609];
                
                r_data[28611] <= r_data[28610];
                
                r_data[28612] <= r_data[28611];
                
                r_data[28613] <= r_data[28612];
                
                r_data[28614] <= r_data[28613];
                
                r_data[28615] <= r_data[28614];
                
                r_data[28616] <= r_data[28615];
                
                r_data[28617] <= r_data[28616];
                
                r_data[28618] <= r_data[28617];
                
                r_data[28619] <= r_data[28618];
                
                r_data[28620] <= r_data[28619];
                
                r_data[28621] <= r_data[28620];
                
                r_data[28622] <= r_data[28621];
                
                r_data[28623] <= r_data[28622];
                
                r_data[28624] <= r_data[28623];
                
                r_data[28625] <= r_data[28624];
                
                r_data[28626] <= r_data[28625];
                
                r_data[28627] <= r_data[28626];
                
                r_data[28628] <= r_data[28627];
                
                r_data[28629] <= r_data[28628];
                
                r_data[28630] <= r_data[28629];
                
                r_data[28631] <= r_data[28630];
                
                r_data[28632] <= r_data[28631];
                
                r_data[28633] <= r_data[28632];
                
                r_data[28634] <= r_data[28633];
                
                r_data[28635] <= r_data[28634];
                
                r_data[28636] <= r_data[28635];
                
                r_data[28637] <= r_data[28636];
                
                r_data[28638] <= r_data[28637];
                
                r_data[28639] <= r_data[28638];
                
                r_data[28640] <= r_data[28639];
                
                r_data[28641] <= r_data[28640];
                
                r_data[28642] <= r_data[28641];
                
                r_data[28643] <= r_data[28642];
                
                r_data[28644] <= r_data[28643];
                
                r_data[28645] <= r_data[28644];
                
                r_data[28646] <= r_data[28645];
                
                r_data[28647] <= r_data[28646];
                
                r_data[28648] <= r_data[28647];
                
                r_data[28649] <= r_data[28648];
                
                r_data[28650] <= r_data[28649];
                
                r_data[28651] <= r_data[28650];
                
                r_data[28652] <= r_data[28651];
                
                r_data[28653] <= r_data[28652];
                
                r_data[28654] <= r_data[28653];
                
                r_data[28655] <= r_data[28654];
                
                r_data[28656] <= r_data[28655];
                
                r_data[28657] <= r_data[28656];
                
                r_data[28658] <= r_data[28657];
                
                r_data[28659] <= r_data[28658];
                
                r_data[28660] <= r_data[28659];
                
                r_data[28661] <= r_data[28660];
                
                r_data[28662] <= r_data[28661];
                
                r_data[28663] <= r_data[28662];
                
                r_data[28664] <= r_data[28663];
                
                r_data[28665] <= r_data[28664];
                
                r_data[28666] <= r_data[28665];
                
                r_data[28667] <= r_data[28666];
                
                r_data[28668] <= r_data[28667];
                
                r_data[28669] <= r_data[28668];
                
                r_data[28670] <= r_data[28669];
                
                r_data[28671] <= r_data[28670];
                
                r_data[28672] <= r_data[28671];
                
                r_data[28673] <= r_data[28672];
                
                r_data[28674] <= r_data[28673];
                
                r_data[28675] <= r_data[28674];
                
                r_data[28676] <= r_data[28675];
                
                r_data[28677] <= r_data[28676];
                
                r_data[28678] <= r_data[28677];
                
                r_data[28679] <= r_data[28678];
                
                r_data[28680] <= r_data[28679];
                
                r_data[28681] <= r_data[28680];
                
                r_data[28682] <= r_data[28681];
                
                r_data[28683] <= r_data[28682];
                
                r_data[28684] <= r_data[28683];
                
                r_data[28685] <= r_data[28684];
                
                r_data[28686] <= r_data[28685];
                
                r_data[28687] <= r_data[28686];
                
                r_data[28688] <= r_data[28687];
                
                r_data[28689] <= r_data[28688];
                
                r_data[28690] <= r_data[28689];
                
                r_data[28691] <= r_data[28690];
                
                r_data[28692] <= r_data[28691];
                
                r_data[28693] <= r_data[28692];
                
                r_data[28694] <= r_data[28693];
                
                r_data[28695] <= r_data[28694];
                
                r_data[28696] <= r_data[28695];
                
                r_data[28697] <= r_data[28696];
                
                r_data[28698] <= r_data[28697];
                
                r_data[28699] <= r_data[28698];
                
                r_data[28700] <= r_data[28699];
                
                r_data[28701] <= r_data[28700];
                
                r_data[28702] <= r_data[28701];
                
                r_data[28703] <= r_data[28702];
                
                r_data[28704] <= r_data[28703];
                
                r_data[28705] <= r_data[28704];
                
                r_data[28706] <= r_data[28705];
                
                r_data[28707] <= r_data[28706];
                
                r_data[28708] <= r_data[28707];
                
                r_data[28709] <= r_data[28708];
                
                r_data[28710] <= r_data[28709];
                
                r_data[28711] <= r_data[28710];
                
                r_data[28712] <= r_data[28711];
                
                r_data[28713] <= r_data[28712];
                
                r_data[28714] <= r_data[28713];
                
                r_data[28715] <= r_data[28714];
                
                r_data[28716] <= r_data[28715];
                
                r_data[28717] <= r_data[28716];
                
                r_data[28718] <= r_data[28717];
                
                r_data[28719] <= r_data[28718];
                
                r_data[28720] <= r_data[28719];
                
                r_data[28721] <= r_data[28720];
                
                r_data[28722] <= r_data[28721];
                
                r_data[28723] <= r_data[28722];
                
                r_data[28724] <= r_data[28723];
                
                r_data[28725] <= r_data[28724];
                
                r_data[28726] <= r_data[28725];
                
                r_data[28727] <= r_data[28726];
                
                r_data[28728] <= r_data[28727];
                
                r_data[28729] <= r_data[28728];
                
                r_data[28730] <= r_data[28729];
                
                r_data[28731] <= r_data[28730];
                
                r_data[28732] <= r_data[28731];
                
                r_data[28733] <= r_data[28732];
                
                r_data[28734] <= r_data[28733];
                
                r_data[28735] <= r_data[28734];
                
                r_data[28736] <= r_data[28735];
                
                r_data[28737] <= r_data[28736];
                
                r_data[28738] <= r_data[28737];
                
                r_data[28739] <= r_data[28738];
                
                r_data[28740] <= r_data[28739];
                
                r_data[28741] <= r_data[28740];
                
                r_data[28742] <= r_data[28741];
                
                r_data[28743] <= r_data[28742];
                
                r_data[28744] <= r_data[28743];
                
                r_data[28745] <= r_data[28744];
                
                r_data[28746] <= r_data[28745];
                
                r_data[28747] <= r_data[28746];
                
                r_data[28748] <= r_data[28747];
                
                r_data[28749] <= r_data[28748];
                
                r_data[28750] <= r_data[28749];
                
                r_data[28751] <= r_data[28750];
                
                r_data[28752] <= r_data[28751];
                
                r_data[28753] <= r_data[28752];
                
                r_data[28754] <= r_data[28753];
                
                r_data[28755] <= r_data[28754];
                
                r_data[28756] <= r_data[28755];
                
                r_data[28757] <= r_data[28756];
                
                r_data[28758] <= r_data[28757];
                
                r_data[28759] <= r_data[28758];
                
                r_data[28760] <= r_data[28759];
                
                r_data[28761] <= r_data[28760];
                
                r_data[28762] <= r_data[28761];
                
                r_data[28763] <= r_data[28762];
                
                r_data[28764] <= r_data[28763];
                
                r_data[28765] <= r_data[28764];
                
                r_data[28766] <= r_data[28765];
                
                r_data[28767] <= r_data[28766];
                
                r_data[28768] <= r_data[28767];
                
                r_data[28769] <= r_data[28768];
                
                r_data[28770] <= r_data[28769];
                
                r_data[28771] <= r_data[28770];
                
                r_data[28772] <= r_data[28771];
                
                r_data[28773] <= r_data[28772];
                
                r_data[28774] <= r_data[28773];
                
                r_data[28775] <= r_data[28774];
                
                r_data[28776] <= r_data[28775];
                
                r_data[28777] <= r_data[28776];
                
                r_data[28778] <= r_data[28777];
                
                r_data[28779] <= r_data[28778];
                
                r_data[28780] <= r_data[28779];
                
                r_data[28781] <= r_data[28780];
                
                r_data[28782] <= r_data[28781];
                
                r_data[28783] <= r_data[28782];
                
                r_data[28784] <= r_data[28783];
                
                r_data[28785] <= r_data[28784];
                
                r_data[28786] <= r_data[28785];
                
                r_data[28787] <= r_data[28786];
                
                r_data[28788] <= r_data[28787];
                
                r_data[28789] <= r_data[28788];
                
                r_data[28790] <= r_data[28789];
                
                r_data[28791] <= r_data[28790];
                
                r_data[28792] <= r_data[28791];
                
                r_data[28793] <= r_data[28792];
                
                r_data[28794] <= r_data[28793];
                
                r_data[28795] <= r_data[28794];
                
                r_data[28796] <= r_data[28795];
                
                r_data[28797] <= r_data[28796];
                
                r_data[28798] <= r_data[28797];
                
                r_data[28799] <= r_data[28798];
                
                r_data[28800] <= r_data[28799];
                
                r_data[28801] <= r_data[28800];
                
                r_data[28802] <= r_data[28801];
                
                r_data[28803] <= r_data[28802];
                
                r_data[28804] <= r_data[28803];
                
                r_data[28805] <= r_data[28804];
                
                r_data[28806] <= r_data[28805];
                
                r_data[28807] <= r_data[28806];
                
                r_data[28808] <= r_data[28807];
                
                r_data[28809] <= r_data[28808];
                
                r_data[28810] <= r_data[28809];
                
                r_data[28811] <= r_data[28810];
                
                r_data[28812] <= r_data[28811];
                
                r_data[28813] <= r_data[28812];
                
                r_data[28814] <= r_data[28813];
                
                r_data[28815] <= r_data[28814];
                
                r_data[28816] <= r_data[28815];
                
                r_data[28817] <= r_data[28816];
                
                r_data[28818] <= r_data[28817];
                
                r_data[28819] <= r_data[28818];
                
                r_data[28820] <= r_data[28819];
                
                r_data[28821] <= r_data[28820];
                
                r_data[28822] <= r_data[28821];
                
                r_data[28823] <= r_data[28822];
                
                r_data[28824] <= r_data[28823];
                
                r_data[28825] <= r_data[28824];
                
                r_data[28826] <= r_data[28825];
                
                r_data[28827] <= r_data[28826];
                
                r_data[28828] <= r_data[28827];
                
                r_data[28829] <= r_data[28828];
                
                r_data[28830] <= r_data[28829];
                
                r_data[28831] <= r_data[28830];
                
                r_data[28832] <= r_data[28831];
                
                r_data[28833] <= r_data[28832];
                
                r_data[28834] <= r_data[28833];
                
                r_data[28835] <= r_data[28834];
                
                r_data[28836] <= r_data[28835];
                
                r_data[28837] <= r_data[28836];
                
                r_data[28838] <= r_data[28837];
                
                r_data[28839] <= r_data[28838];
                
                r_data[28840] <= r_data[28839];
                
                r_data[28841] <= r_data[28840];
                
                r_data[28842] <= r_data[28841];
                
                r_data[28843] <= r_data[28842];
                
                r_data[28844] <= r_data[28843];
                
                r_data[28845] <= r_data[28844];
                
                r_data[28846] <= r_data[28845];
                
                r_data[28847] <= r_data[28846];
                
                r_data[28848] <= r_data[28847];
                
                r_data[28849] <= r_data[28848];
                
                r_data[28850] <= r_data[28849];
                
                r_data[28851] <= r_data[28850];
                
                r_data[28852] <= r_data[28851];
                
                r_data[28853] <= r_data[28852];
                
                r_data[28854] <= r_data[28853];
                
                r_data[28855] <= r_data[28854];
                
                r_data[28856] <= r_data[28855];
                
                r_data[28857] <= r_data[28856];
                
                r_data[28858] <= r_data[28857];
                
                r_data[28859] <= r_data[28858];
                
                r_data[28860] <= r_data[28859];
                
                r_data[28861] <= r_data[28860];
                
                r_data[28862] <= r_data[28861];
                
                r_data[28863] <= r_data[28862];
                
                r_data[28864] <= r_data[28863];
                
                r_data[28865] <= r_data[28864];
                
                r_data[28866] <= r_data[28865];
                
                r_data[28867] <= r_data[28866];
                
                r_data[28868] <= r_data[28867];
                
                r_data[28869] <= r_data[28868];
                
                r_data[28870] <= r_data[28869];
                
                r_data[28871] <= r_data[28870];
                
                r_data[28872] <= r_data[28871];
                
                r_data[28873] <= r_data[28872];
                
                r_data[28874] <= r_data[28873];
                
                r_data[28875] <= r_data[28874];
                
                r_data[28876] <= r_data[28875];
                
                r_data[28877] <= r_data[28876];
                
                r_data[28878] <= r_data[28877];
                
                r_data[28879] <= r_data[28878];
                
                r_data[28880] <= r_data[28879];
                
                r_data[28881] <= r_data[28880];
                
                r_data[28882] <= r_data[28881];
                
                r_data[28883] <= r_data[28882];
                
                r_data[28884] <= r_data[28883];
                
                r_data[28885] <= r_data[28884];
                
                r_data[28886] <= r_data[28885];
                
                r_data[28887] <= r_data[28886];
                
                r_data[28888] <= r_data[28887];
                
                r_data[28889] <= r_data[28888];
                
                r_data[28890] <= r_data[28889];
                
                r_data[28891] <= r_data[28890];
                
                r_data[28892] <= r_data[28891];
                
                r_data[28893] <= r_data[28892];
                
                r_data[28894] <= r_data[28893];
                
                r_data[28895] <= r_data[28894];
                
                r_data[28896] <= r_data[28895];
                
                r_data[28897] <= r_data[28896];
                
                r_data[28898] <= r_data[28897];
                
                r_data[28899] <= r_data[28898];
                
                r_data[28900] <= r_data[28899];
                
                r_data[28901] <= r_data[28900];
                
                r_data[28902] <= r_data[28901];
                
                r_data[28903] <= r_data[28902];
                
                r_data[28904] <= r_data[28903];
                
                r_data[28905] <= r_data[28904];
                
                r_data[28906] <= r_data[28905];
                
                r_data[28907] <= r_data[28906];
                
                r_data[28908] <= r_data[28907];
                
                r_data[28909] <= r_data[28908];
                
                r_data[28910] <= r_data[28909];
                
                r_data[28911] <= r_data[28910];
                
                r_data[28912] <= r_data[28911];
                
                r_data[28913] <= r_data[28912];
                
                r_data[28914] <= r_data[28913];
                
                r_data[28915] <= r_data[28914];
                
                r_data[28916] <= r_data[28915];
                
                r_data[28917] <= r_data[28916];
                
                r_data[28918] <= r_data[28917];
                
                r_data[28919] <= r_data[28918];
                
                r_data[28920] <= r_data[28919];
                
                r_data[28921] <= r_data[28920];
                
                r_data[28922] <= r_data[28921];
                
                r_data[28923] <= r_data[28922];
                
                r_data[28924] <= r_data[28923];
                
                r_data[28925] <= r_data[28924];
                
                r_data[28926] <= r_data[28925];
                
                r_data[28927] <= r_data[28926];
                
                r_data[28928] <= r_data[28927];
                
                r_data[28929] <= r_data[28928];
                
                r_data[28930] <= r_data[28929];
                
                r_data[28931] <= r_data[28930];
                
                r_data[28932] <= r_data[28931];
                
                r_data[28933] <= r_data[28932];
                
                r_data[28934] <= r_data[28933];
                
                r_data[28935] <= r_data[28934];
                
                r_data[28936] <= r_data[28935];
                
                r_data[28937] <= r_data[28936];
                
                r_data[28938] <= r_data[28937];
                
                r_data[28939] <= r_data[28938];
                
                r_data[28940] <= r_data[28939];
                
                r_data[28941] <= r_data[28940];
                
                r_data[28942] <= r_data[28941];
                
                r_data[28943] <= r_data[28942];
                
                r_data[28944] <= r_data[28943];
                
                r_data[28945] <= r_data[28944];
                
                r_data[28946] <= r_data[28945];
                
                r_data[28947] <= r_data[28946];
                
                r_data[28948] <= r_data[28947];
                
                r_data[28949] <= r_data[28948];
                
                r_data[28950] <= r_data[28949];
                
                r_data[28951] <= r_data[28950];
                
                r_data[28952] <= r_data[28951];
                
                r_data[28953] <= r_data[28952];
                
                r_data[28954] <= r_data[28953];
                
                r_data[28955] <= r_data[28954];
                
                r_data[28956] <= r_data[28955];
                
                r_data[28957] <= r_data[28956];
                
                r_data[28958] <= r_data[28957];
                
                r_data[28959] <= r_data[28958];
                
                r_data[28960] <= r_data[28959];
                
                r_data[28961] <= r_data[28960];
                
                r_data[28962] <= r_data[28961];
                
                r_data[28963] <= r_data[28962];
                
                r_data[28964] <= r_data[28963];
                
                r_data[28965] <= r_data[28964];
                
                r_data[28966] <= r_data[28965];
                
                r_data[28967] <= r_data[28966];
                
                r_data[28968] <= r_data[28967];
                
                r_data[28969] <= r_data[28968];
                
                r_data[28970] <= r_data[28969];
                
                r_data[28971] <= r_data[28970];
                
                r_data[28972] <= r_data[28971];
                
                r_data[28973] <= r_data[28972];
                
                r_data[28974] <= r_data[28973];
                
                r_data[28975] <= r_data[28974];
                
                r_data[28976] <= r_data[28975];
                
                r_data[28977] <= r_data[28976];
                
                r_data[28978] <= r_data[28977];
                
                r_data[28979] <= r_data[28978];
                
                r_data[28980] <= r_data[28979];
                
                r_data[28981] <= r_data[28980];
                
                r_data[28982] <= r_data[28981];
                
                r_data[28983] <= r_data[28982];
                
                r_data[28984] <= r_data[28983];
                
                r_data[28985] <= r_data[28984];
                
                r_data[28986] <= r_data[28985];
                
                r_data[28987] <= r_data[28986];
                
                r_data[28988] <= r_data[28987];
                
                r_data[28989] <= r_data[28988];
                
                r_data[28990] <= r_data[28989];
                
                r_data[28991] <= r_data[28990];
                
                r_data[28992] <= r_data[28991];
                
                r_data[28993] <= r_data[28992];
                
                r_data[28994] <= r_data[28993];
                
                r_data[28995] <= r_data[28994];
                
                r_data[28996] <= r_data[28995];
                
                r_data[28997] <= r_data[28996];
                
                r_data[28998] <= r_data[28997];
                
                r_data[28999] <= r_data[28998];
                
                r_data[29000] <= r_data[28999];
                
                r_data[29001] <= r_data[29000];
                
                r_data[29002] <= r_data[29001];
                
                r_data[29003] <= r_data[29002];
                
                r_data[29004] <= r_data[29003];
                
                r_data[29005] <= r_data[29004];
                
                r_data[29006] <= r_data[29005];
                
                r_data[29007] <= r_data[29006];
                
                r_data[29008] <= r_data[29007];
                
                r_data[29009] <= r_data[29008];
                
                r_data[29010] <= r_data[29009];
                
                r_data[29011] <= r_data[29010];
                
                r_data[29012] <= r_data[29011];
                
                r_data[29013] <= r_data[29012];
                
                r_data[29014] <= r_data[29013];
                
                r_data[29015] <= r_data[29014];
                
                r_data[29016] <= r_data[29015];
                
                r_data[29017] <= r_data[29016];
                
                r_data[29018] <= r_data[29017];
                
                r_data[29019] <= r_data[29018];
                
                r_data[29020] <= r_data[29019];
                
                r_data[29021] <= r_data[29020];
                
                r_data[29022] <= r_data[29021];
                
                r_data[29023] <= r_data[29022];
                
                r_data[29024] <= r_data[29023];
                
                r_data[29025] <= r_data[29024];
                
                r_data[29026] <= r_data[29025];
                
                r_data[29027] <= r_data[29026];
                
                r_data[29028] <= r_data[29027];
                
                r_data[29029] <= r_data[29028];
                
                r_data[29030] <= r_data[29029];
                
                r_data[29031] <= r_data[29030];
                
                r_data[29032] <= r_data[29031];
                
                r_data[29033] <= r_data[29032];
                
                r_data[29034] <= r_data[29033];
                
                r_data[29035] <= r_data[29034];
                
                r_data[29036] <= r_data[29035];
                
                r_data[29037] <= r_data[29036];
                
                r_data[29038] <= r_data[29037];
                
                r_data[29039] <= r_data[29038];
                
                r_data[29040] <= r_data[29039];
                
                r_data[29041] <= r_data[29040];
                
                r_data[29042] <= r_data[29041];
                
                r_data[29043] <= r_data[29042];
                
                r_data[29044] <= r_data[29043];
                
                r_data[29045] <= r_data[29044];
                
                r_data[29046] <= r_data[29045];
                
                r_data[29047] <= r_data[29046];
                
                r_data[29048] <= r_data[29047];
                
                r_data[29049] <= r_data[29048];
                
                r_data[29050] <= r_data[29049];
                
                r_data[29051] <= r_data[29050];
                
                r_data[29052] <= r_data[29051];
                
                r_data[29053] <= r_data[29052];
                
                r_data[29054] <= r_data[29053];
                
                r_data[29055] <= r_data[29054];
                
                r_data[29056] <= r_data[29055];
                
                r_data[29057] <= r_data[29056];
                
                r_data[29058] <= r_data[29057];
                
                r_data[29059] <= r_data[29058];
                
                r_data[29060] <= r_data[29059];
                
                r_data[29061] <= r_data[29060];
                
                r_data[29062] <= r_data[29061];
                
                r_data[29063] <= r_data[29062];
                
                r_data[29064] <= r_data[29063];
                
                r_data[29065] <= r_data[29064];
                
                r_data[29066] <= r_data[29065];
                
                r_data[29067] <= r_data[29066];
                
                r_data[29068] <= r_data[29067];
                
                r_data[29069] <= r_data[29068];
                
                r_data[29070] <= r_data[29069];
                
                r_data[29071] <= r_data[29070];
                
                r_data[29072] <= r_data[29071];
                
                r_data[29073] <= r_data[29072];
                
                r_data[29074] <= r_data[29073];
                
                r_data[29075] <= r_data[29074];
                
                r_data[29076] <= r_data[29075];
                
                r_data[29077] <= r_data[29076];
                
                r_data[29078] <= r_data[29077];
                
                r_data[29079] <= r_data[29078];
                
                r_data[29080] <= r_data[29079];
                
                r_data[29081] <= r_data[29080];
                
                r_data[29082] <= r_data[29081];
                
                r_data[29083] <= r_data[29082];
                
                r_data[29084] <= r_data[29083];
                
                r_data[29085] <= r_data[29084];
                
                r_data[29086] <= r_data[29085];
                
                r_data[29087] <= r_data[29086];
                
                r_data[29088] <= r_data[29087];
                
                r_data[29089] <= r_data[29088];
                
                r_data[29090] <= r_data[29089];
                
                r_data[29091] <= r_data[29090];
                
                r_data[29092] <= r_data[29091];
                
                r_data[29093] <= r_data[29092];
                
                r_data[29094] <= r_data[29093];
                
                r_data[29095] <= r_data[29094];
                
                r_data[29096] <= r_data[29095];
                
                r_data[29097] <= r_data[29096];
                
                r_data[29098] <= r_data[29097];
                
                r_data[29099] <= r_data[29098];
                
                r_data[29100] <= r_data[29099];
                
                r_data[29101] <= r_data[29100];
                
                r_data[29102] <= r_data[29101];
                
                r_data[29103] <= r_data[29102];
                
                r_data[29104] <= r_data[29103];
                
                r_data[29105] <= r_data[29104];
                
                r_data[29106] <= r_data[29105];
                
                r_data[29107] <= r_data[29106];
                
                r_data[29108] <= r_data[29107];
                
                r_data[29109] <= r_data[29108];
                
                r_data[29110] <= r_data[29109];
                
                r_data[29111] <= r_data[29110];
                
                r_data[29112] <= r_data[29111];
                
                r_data[29113] <= r_data[29112];
                
                r_data[29114] <= r_data[29113];
                
                r_data[29115] <= r_data[29114];
                
                r_data[29116] <= r_data[29115];
                
                r_data[29117] <= r_data[29116];
                
                r_data[29118] <= r_data[29117];
                
                r_data[29119] <= r_data[29118];
                
                r_data[29120] <= r_data[29119];
                
                r_data[29121] <= r_data[29120];
                
                r_data[29122] <= r_data[29121];
                
                r_data[29123] <= r_data[29122];
                
                r_data[29124] <= r_data[29123];
                
                r_data[29125] <= r_data[29124];
                
                r_data[29126] <= r_data[29125];
                
                r_data[29127] <= r_data[29126];
                
                r_data[29128] <= r_data[29127];
                
                r_data[29129] <= r_data[29128];
                
                r_data[29130] <= r_data[29129];
                
                r_data[29131] <= r_data[29130];
                
                r_data[29132] <= r_data[29131];
                
                r_data[29133] <= r_data[29132];
                
                r_data[29134] <= r_data[29133];
                
                r_data[29135] <= r_data[29134];
                
                r_data[29136] <= r_data[29135];
                
                r_data[29137] <= r_data[29136];
                
                r_data[29138] <= r_data[29137];
                
                r_data[29139] <= r_data[29138];
                
                r_data[29140] <= r_data[29139];
                
                r_data[29141] <= r_data[29140];
                
                r_data[29142] <= r_data[29141];
                
                r_data[29143] <= r_data[29142];
                
                r_data[29144] <= r_data[29143];
                
                r_data[29145] <= r_data[29144];
                
                r_data[29146] <= r_data[29145];
                
                r_data[29147] <= r_data[29146];
                
                r_data[29148] <= r_data[29147];
                
                r_data[29149] <= r_data[29148];
                
                r_data[29150] <= r_data[29149];
                
                r_data[29151] <= r_data[29150];
                
                r_data[29152] <= r_data[29151];
                
                r_data[29153] <= r_data[29152];
                
                r_data[29154] <= r_data[29153];
                
                r_data[29155] <= r_data[29154];
                
                r_data[29156] <= r_data[29155];
                
                r_data[29157] <= r_data[29156];
                
                r_data[29158] <= r_data[29157];
                
                r_data[29159] <= r_data[29158];
                
                r_data[29160] <= r_data[29159];
                
                r_data[29161] <= r_data[29160];
                
                r_data[29162] <= r_data[29161];
                
                r_data[29163] <= r_data[29162];
                
                r_data[29164] <= r_data[29163];
                
                r_data[29165] <= r_data[29164];
                
                r_data[29166] <= r_data[29165];
                
                r_data[29167] <= r_data[29166];
                
                r_data[29168] <= r_data[29167];
                
                r_data[29169] <= r_data[29168];
                
                r_data[29170] <= r_data[29169];
                
                r_data[29171] <= r_data[29170];
                
                r_data[29172] <= r_data[29171];
                
                r_data[29173] <= r_data[29172];
                
                r_data[29174] <= r_data[29173];
                
                r_data[29175] <= r_data[29174];
                
                r_data[29176] <= r_data[29175];
                
                r_data[29177] <= r_data[29176];
                
                r_data[29178] <= r_data[29177];
                
                r_data[29179] <= r_data[29178];
                
                r_data[29180] <= r_data[29179];
                
                r_data[29181] <= r_data[29180];
                
                r_data[29182] <= r_data[29181];
                
                r_data[29183] <= r_data[29182];
                
                r_data[29184] <= r_data[29183];
                
                r_data[29185] <= r_data[29184];
                
                r_data[29186] <= r_data[29185];
                
                r_data[29187] <= r_data[29186];
                
                r_data[29188] <= r_data[29187];
                
                r_data[29189] <= r_data[29188];
                
                r_data[29190] <= r_data[29189];
                
                r_data[29191] <= r_data[29190];
                
                r_data[29192] <= r_data[29191];
                
                r_data[29193] <= r_data[29192];
                
                r_data[29194] <= r_data[29193];
                
                r_data[29195] <= r_data[29194];
                
                r_data[29196] <= r_data[29195];
                
                r_data[29197] <= r_data[29196];
                
                r_data[29198] <= r_data[29197];
                
                r_data[29199] <= r_data[29198];
                
                r_data[29200] <= r_data[29199];
                
                r_data[29201] <= r_data[29200];
                
                r_data[29202] <= r_data[29201];
                
                r_data[29203] <= r_data[29202];
                
                r_data[29204] <= r_data[29203];
                
                r_data[29205] <= r_data[29204];
                
                r_data[29206] <= r_data[29205];
                
                r_data[29207] <= r_data[29206];
                
                r_data[29208] <= r_data[29207];
                
                r_data[29209] <= r_data[29208];
                
                r_data[29210] <= r_data[29209];
                
                r_data[29211] <= r_data[29210];
                
                r_data[29212] <= r_data[29211];
                
                r_data[29213] <= r_data[29212];
                
                r_data[29214] <= r_data[29213];
                
                r_data[29215] <= r_data[29214];
                
                r_data[29216] <= r_data[29215];
                
                r_data[29217] <= r_data[29216];
                
                r_data[29218] <= r_data[29217];
                
                r_data[29219] <= r_data[29218];
                
                r_data[29220] <= r_data[29219];
                
                r_data[29221] <= r_data[29220];
                
                r_data[29222] <= r_data[29221];
                
                r_data[29223] <= r_data[29222];
                
                r_data[29224] <= r_data[29223];
                
                r_data[29225] <= r_data[29224];
                
                r_data[29226] <= r_data[29225];
                
                r_data[29227] <= r_data[29226];
                
                r_data[29228] <= r_data[29227];
                
                r_data[29229] <= r_data[29228];
                
                r_data[29230] <= r_data[29229];
                
                r_data[29231] <= r_data[29230];
                
                r_data[29232] <= r_data[29231];
                
                r_data[29233] <= r_data[29232];
                
                r_data[29234] <= r_data[29233];
                
                r_data[29235] <= r_data[29234];
                
                r_data[29236] <= r_data[29235];
                
                r_data[29237] <= r_data[29236];
                
                r_data[29238] <= r_data[29237];
                
                r_data[29239] <= r_data[29238];
                
                r_data[29240] <= r_data[29239];
                
                r_data[29241] <= r_data[29240];
                
                r_data[29242] <= r_data[29241];
                
                r_data[29243] <= r_data[29242];
                
                r_data[29244] <= r_data[29243];
                
                r_data[29245] <= r_data[29244];
                
                r_data[29246] <= r_data[29245];
                
                r_data[29247] <= r_data[29246];
                
                r_data[29248] <= r_data[29247];
                
                r_data[29249] <= r_data[29248];
                
                r_data[29250] <= r_data[29249];
                
                r_data[29251] <= r_data[29250];
                
                r_data[29252] <= r_data[29251];
                
                r_data[29253] <= r_data[29252];
                
                r_data[29254] <= r_data[29253];
                
                r_data[29255] <= r_data[29254];
                
                r_data[29256] <= r_data[29255];
                
                r_data[29257] <= r_data[29256];
                
                r_data[29258] <= r_data[29257];
                
                r_data[29259] <= r_data[29258];
                
                r_data[29260] <= r_data[29259];
                
                r_data[29261] <= r_data[29260];
                
                r_data[29262] <= r_data[29261];
                
                r_data[29263] <= r_data[29262];
                
                r_data[29264] <= r_data[29263];
                
                r_data[29265] <= r_data[29264];
                
                r_data[29266] <= r_data[29265];
                
                r_data[29267] <= r_data[29266];
                
                r_data[29268] <= r_data[29267];
                
                r_data[29269] <= r_data[29268];
                
                r_data[29270] <= r_data[29269];
                
                r_data[29271] <= r_data[29270];
                
                r_data[29272] <= r_data[29271];
                
                r_data[29273] <= r_data[29272];
                
                r_data[29274] <= r_data[29273];
                
                r_data[29275] <= r_data[29274];
                
                r_data[29276] <= r_data[29275];
                
                r_data[29277] <= r_data[29276];
                
                r_data[29278] <= r_data[29277];
                
                r_data[29279] <= r_data[29278];
                
                r_data[29280] <= r_data[29279];
                
                r_data[29281] <= r_data[29280];
                
                r_data[29282] <= r_data[29281];
                
                r_data[29283] <= r_data[29282];
                
                r_data[29284] <= r_data[29283];
                
                r_data[29285] <= r_data[29284];
                
                r_data[29286] <= r_data[29285];
                
                r_data[29287] <= r_data[29286];
                
                r_data[29288] <= r_data[29287];
                
                r_data[29289] <= r_data[29288];
                
                r_data[29290] <= r_data[29289];
                
                r_data[29291] <= r_data[29290];
                
                r_data[29292] <= r_data[29291];
                
                r_data[29293] <= r_data[29292];
                
                r_data[29294] <= r_data[29293];
                
                r_data[29295] <= r_data[29294];
                
                r_data[29296] <= r_data[29295];
                
                r_data[29297] <= r_data[29296];
                
                r_data[29298] <= r_data[29297];
                
                r_data[29299] <= r_data[29298];
                
                r_data[29300] <= r_data[29299];
                
                r_data[29301] <= r_data[29300];
                
                r_data[29302] <= r_data[29301];
                
                r_data[29303] <= r_data[29302];
                
                r_data[29304] <= r_data[29303];
                
                r_data[29305] <= r_data[29304];
                
                r_data[29306] <= r_data[29305];
                
                r_data[29307] <= r_data[29306];
                
                r_data[29308] <= r_data[29307];
                
                r_data[29309] <= r_data[29308];
                
                r_data[29310] <= r_data[29309];
                
                r_data[29311] <= r_data[29310];
                
                r_data[29312] <= r_data[29311];
                
                r_data[29313] <= r_data[29312];
                
                r_data[29314] <= r_data[29313];
                
                r_data[29315] <= r_data[29314];
                
                r_data[29316] <= r_data[29315];
                
                r_data[29317] <= r_data[29316];
                
                r_data[29318] <= r_data[29317];
                
                r_data[29319] <= r_data[29318];
                
                r_data[29320] <= r_data[29319];
                
                r_data[29321] <= r_data[29320];
                
                r_data[29322] <= r_data[29321];
                
                r_data[29323] <= r_data[29322];
                
                r_data[29324] <= r_data[29323];
                
                r_data[29325] <= r_data[29324];
                
                r_data[29326] <= r_data[29325];
                
                r_data[29327] <= r_data[29326];
                
                r_data[29328] <= r_data[29327];
                
                r_data[29329] <= r_data[29328];
                
                r_data[29330] <= r_data[29329];
                
                r_data[29331] <= r_data[29330];
                
                r_data[29332] <= r_data[29331];
                
                r_data[29333] <= r_data[29332];
                
                r_data[29334] <= r_data[29333];
                
                r_data[29335] <= r_data[29334];
                
                r_data[29336] <= r_data[29335];
                
                r_data[29337] <= r_data[29336];
                
                r_data[29338] <= r_data[29337];
                
                r_data[29339] <= r_data[29338];
                
                r_data[29340] <= r_data[29339];
                
                r_data[29341] <= r_data[29340];
                
                r_data[29342] <= r_data[29341];
                
                r_data[29343] <= r_data[29342];
                
                r_data[29344] <= r_data[29343];
                
                r_data[29345] <= r_data[29344];
                
                r_data[29346] <= r_data[29345];
                
                r_data[29347] <= r_data[29346];
                
                r_data[29348] <= r_data[29347];
                
                r_data[29349] <= r_data[29348];
                
                r_data[29350] <= r_data[29349];
                
                r_data[29351] <= r_data[29350];
                
                r_data[29352] <= r_data[29351];
                
                r_data[29353] <= r_data[29352];
                
                r_data[29354] <= r_data[29353];
                
                r_data[29355] <= r_data[29354];
                
                r_data[29356] <= r_data[29355];
                
                r_data[29357] <= r_data[29356];
                
                r_data[29358] <= r_data[29357];
                
                r_data[29359] <= r_data[29358];
                
                r_data[29360] <= r_data[29359];
                
                r_data[29361] <= r_data[29360];
                
                r_data[29362] <= r_data[29361];
                
                r_data[29363] <= r_data[29362];
                
                r_data[29364] <= r_data[29363];
                
                r_data[29365] <= r_data[29364];
                
                r_data[29366] <= r_data[29365];
                
                r_data[29367] <= r_data[29366];
                
                r_data[29368] <= r_data[29367];
                
                r_data[29369] <= r_data[29368];
                
                r_data[29370] <= r_data[29369];
                
                r_data[29371] <= r_data[29370];
                
                r_data[29372] <= r_data[29371];
                
                r_data[29373] <= r_data[29372];
                
                r_data[29374] <= r_data[29373];
                
                r_data[29375] <= r_data[29374];
                
                r_data[29376] <= r_data[29375];
                
                r_data[29377] <= r_data[29376];
                
                r_data[29378] <= r_data[29377];
                
                r_data[29379] <= r_data[29378];
                
                r_data[29380] <= r_data[29379];
                
                r_data[29381] <= r_data[29380];
                
                r_data[29382] <= r_data[29381];
                
                r_data[29383] <= r_data[29382];
                
                r_data[29384] <= r_data[29383];
                
                r_data[29385] <= r_data[29384];
                
                r_data[29386] <= r_data[29385];
                
                r_data[29387] <= r_data[29386];
                
                r_data[29388] <= r_data[29387];
                
                r_data[29389] <= r_data[29388];
                
                r_data[29390] <= r_data[29389];
                
                r_data[29391] <= r_data[29390];
                
                r_data[29392] <= r_data[29391];
                
                r_data[29393] <= r_data[29392];
                
                r_data[29394] <= r_data[29393];
                
                r_data[29395] <= r_data[29394];
                
                r_data[29396] <= r_data[29395];
                
                r_data[29397] <= r_data[29396];
                
                r_data[29398] <= r_data[29397];
                
                r_data[29399] <= r_data[29398];
                
                r_data[29400] <= r_data[29399];
                
                r_data[29401] <= r_data[29400];
                
                r_data[29402] <= r_data[29401];
                
                r_data[29403] <= r_data[29402];
                
                r_data[29404] <= r_data[29403];
                
                r_data[29405] <= r_data[29404];
                
                r_data[29406] <= r_data[29405];
                
                r_data[29407] <= r_data[29406];
                
                r_data[29408] <= r_data[29407];
                
                r_data[29409] <= r_data[29408];
                
                r_data[29410] <= r_data[29409];
                
                r_data[29411] <= r_data[29410];
                
                r_data[29412] <= r_data[29411];
                
                r_data[29413] <= r_data[29412];
                
                r_data[29414] <= r_data[29413];
                
                r_data[29415] <= r_data[29414];
                
                r_data[29416] <= r_data[29415];
                
                r_data[29417] <= r_data[29416];
                
                r_data[29418] <= r_data[29417];
                
                r_data[29419] <= r_data[29418];
                
                r_data[29420] <= r_data[29419];
                
                r_data[29421] <= r_data[29420];
                
                r_data[29422] <= r_data[29421];
                
                r_data[29423] <= r_data[29422];
                
                r_data[29424] <= r_data[29423];
                
                r_data[29425] <= r_data[29424];
                
                r_data[29426] <= r_data[29425];
                
                r_data[29427] <= r_data[29426];
                
                r_data[29428] <= r_data[29427];
                
                r_data[29429] <= r_data[29428];
                
                r_data[29430] <= r_data[29429];
                
                r_data[29431] <= r_data[29430];
                
                r_data[29432] <= r_data[29431];
                
                r_data[29433] <= r_data[29432];
                
                r_data[29434] <= r_data[29433];
                
                r_data[29435] <= r_data[29434];
                
                r_data[29436] <= r_data[29435];
                
                r_data[29437] <= r_data[29436];
                
                r_data[29438] <= r_data[29437];
                
                r_data[29439] <= r_data[29438];
                
                r_data[29440] <= r_data[29439];
                
                r_data[29441] <= r_data[29440];
                
                r_data[29442] <= r_data[29441];
                
                r_data[29443] <= r_data[29442];
                
                r_data[29444] <= r_data[29443];
                
                r_data[29445] <= r_data[29444];
                
                r_data[29446] <= r_data[29445];
                
                r_data[29447] <= r_data[29446];
                
                r_data[29448] <= r_data[29447];
                
                r_data[29449] <= r_data[29448];
                
                r_data[29450] <= r_data[29449];
                
                r_data[29451] <= r_data[29450];
                
                r_data[29452] <= r_data[29451];
                
                r_data[29453] <= r_data[29452];
                
                r_data[29454] <= r_data[29453];
                
                r_data[29455] <= r_data[29454];
                
                r_data[29456] <= r_data[29455];
                
                r_data[29457] <= r_data[29456];
                
                r_data[29458] <= r_data[29457];
                
                r_data[29459] <= r_data[29458];
                
                r_data[29460] <= r_data[29459];
                
                r_data[29461] <= r_data[29460];
                
                r_data[29462] <= r_data[29461];
                
                r_data[29463] <= r_data[29462];
                
                r_data[29464] <= r_data[29463];
                
                r_data[29465] <= r_data[29464];
                
                r_data[29466] <= r_data[29465];
                
                r_data[29467] <= r_data[29466];
                
                r_data[29468] <= r_data[29467];
                
                r_data[29469] <= r_data[29468];
                
                r_data[29470] <= r_data[29469];
                
                r_data[29471] <= r_data[29470];
                
                r_data[29472] <= r_data[29471];
                
                r_data[29473] <= r_data[29472];
                
                r_data[29474] <= r_data[29473];
                
                r_data[29475] <= r_data[29474];
                
                r_data[29476] <= r_data[29475];
                
                r_data[29477] <= r_data[29476];
                
                r_data[29478] <= r_data[29477];
                
                r_data[29479] <= r_data[29478];
                
                r_data[29480] <= r_data[29479];
                
                r_data[29481] <= r_data[29480];
                
                r_data[29482] <= r_data[29481];
                
                r_data[29483] <= r_data[29482];
                
                r_data[29484] <= r_data[29483];
                
                r_data[29485] <= r_data[29484];
                
                r_data[29486] <= r_data[29485];
                
                r_data[29487] <= r_data[29486];
                
                r_data[29488] <= r_data[29487];
                
                r_data[29489] <= r_data[29488];
                
                r_data[29490] <= r_data[29489];
                
                r_data[29491] <= r_data[29490];
                
                r_data[29492] <= r_data[29491];
                
                r_data[29493] <= r_data[29492];
                
                r_data[29494] <= r_data[29493];
                
                r_data[29495] <= r_data[29494];
                
                r_data[29496] <= r_data[29495];
                
                r_data[29497] <= r_data[29496];
                
                r_data[29498] <= r_data[29497];
                
                r_data[29499] <= r_data[29498];
                
                r_data[29500] <= r_data[29499];
                
                r_data[29501] <= r_data[29500];
                
                r_data[29502] <= r_data[29501];
                
                r_data[29503] <= r_data[29502];
                
                r_data[29504] <= r_data[29503];
                
                r_data[29505] <= r_data[29504];
                
                r_data[29506] <= r_data[29505];
                
                r_data[29507] <= r_data[29506];
                
                r_data[29508] <= r_data[29507];
                
                r_data[29509] <= r_data[29508];
                
                r_data[29510] <= r_data[29509];
                
                r_data[29511] <= r_data[29510];
                
                r_data[29512] <= r_data[29511];
                
                r_data[29513] <= r_data[29512];
                
                r_data[29514] <= r_data[29513];
                
                r_data[29515] <= r_data[29514];
                
                r_data[29516] <= r_data[29515];
                
                r_data[29517] <= r_data[29516];
                
                r_data[29518] <= r_data[29517];
                
                r_data[29519] <= r_data[29518];
                
                r_data[29520] <= r_data[29519];
                
                r_data[29521] <= r_data[29520];
                
                r_data[29522] <= r_data[29521];
                
                r_data[29523] <= r_data[29522];
                
                r_data[29524] <= r_data[29523];
                
                r_data[29525] <= r_data[29524];
                
                r_data[29526] <= r_data[29525];
                
                r_data[29527] <= r_data[29526];
                
                r_data[29528] <= r_data[29527];
                
                r_data[29529] <= r_data[29528];
                
                r_data[29530] <= r_data[29529];
                
                r_data[29531] <= r_data[29530];
                
                r_data[29532] <= r_data[29531];
                
                r_data[29533] <= r_data[29532];
                
                r_data[29534] <= r_data[29533];
                
                r_data[29535] <= r_data[29534];
                
                r_data[29536] <= r_data[29535];
                
                r_data[29537] <= r_data[29536];
                
                r_data[29538] <= r_data[29537];
                
                r_data[29539] <= r_data[29538];
                
                r_data[29540] <= r_data[29539];
                
                r_data[29541] <= r_data[29540];
                
                r_data[29542] <= r_data[29541];
                
                r_data[29543] <= r_data[29542];
                
                r_data[29544] <= r_data[29543];
                
                r_data[29545] <= r_data[29544];
                
                r_data[29546] <= r_data[29545];
                
                r_data[29547] <= r_data[29546];
                
                r_data[29548] <= r_data[29547];
                
                r_data[29549] <= r_data[29548];
                
                r_data[29550] <= r_data[29549];
                
                r_data[29551] <= r_data[29550];
                
                r_data[29552] <= r_data[29551];
                
                r_data[29553] <= r_data[29552];
                
                r_data[29554] <= r_data[29553];
                
                r_data[29555] <= r_data[29554];
                
                r_data[29556] <= r_data[29555];
                
                r_data[29557] <= r_data[29556];
                
                r_data[29558] <= r_data[29557];
                
                r_data[29559] <= r_data[29558];
                
                r_data[29560] <= r_data[29559];
                
                r_data[29561] <= r_data[29560];
                
                r_data[29562] <= r_data[29561];
                
                r_data[29563] <= r_data[29562];
                
                r_data[29564] <= r_data[29563];
                
                r_data[29565] <= r_data[29564];
                
                r_data[29566] <= r_data[29565];
                
                r_data[29567] <= r_data[29566];
                
                r_data[29568] <= r_data[29567];
                
                r_data[29569] <= r_data[29568];
                
                r_data[29570] <= r_data[29569];
                
                r_data[29571] <= r_data[29570];
                
                r_data[29572] <= r_data[29571];
                
                r_data[29573] <= r_data[29572];
                
                r_data[29574] <= r_data[29573];
                
                r_data[29575] <= r_data[29574];
                
                r_data[29576] <= r_data[29575];
                
                r_data[29577] <= r_data[29576];
                
                r_data[29578] <= r_data[29577];
                
                r_data[29579] <= r_data[29578];
                
                r_data[29580] <= r_data[29579];
                
                r_data[29581] <= r_data[29580];
                
                r_data[29582] <= r_data[29581];
                
                r_data[29583] <= r_data[29582];
                
                r_data[29584] <= r_data[29583];
                
                r_data[29585] <= r_data[29584];
                
                r_data[29586] <= r_data[29585];
                
                r_data[29587] <= r_data[29586];
                
                r_data[29588] <= r_data[29587];
                
                r_data[29589] <= r_data[29588];
                
                r_data[29590] <= r_data[29589];
                
                r_data[29591] <= r_data[29590];
                
                r_data[29592] <= r_data[29591];
                
                r_data[29593] <= r_data[29592];
                
                r_data[29594] <= r_data[29593];
                
                r_data[29595] <= r_data[29594];
                
                r_data[29596] <= r_data[29595];
                
                r_data[29597] <= r_data[29596];
                
                r_data[29598] <= r_data[29597];
                
                r_data[29599] <= r_data[29598];
                
                r_data[29600] <= r_data[29599];
                
                r_data[29601] <= r_data[29600];
                
                r_data[29602] <= r_data[29601];
                
                r_data[29603] <= r_data[29602];
                
                r_data[29604] <= r_data[29603];
                
                r_data[29605] <= r_data[29604];
                
                r_data[29606] <= r_data[29605];
                
                r_data[29607] <= r_data[29606];
                
                r_data[29608] <= r_data[29607];
                
                r_data[29609] <= r_data[29608];
                
                r_data[29610] <= r_data[29609];
                
                r_data[29611] <= r_data[29610];
                
                r_data[29612] <= r_data[29611];
                
                r_data[29613] <= r_data[29612];
                
                r_data[29614] <= r_data[29613];
                
                r_data[29615] <= r_data[29614];
                
                r_data[29616] <= r_data[29615];
                
                r_data[29617] <= r_data[29616];
                
                r_data[29618] <= r_data[29617];
                
                r_data[29619] <= r_data[29618];
                
                r_data[29620] <= r_data[29619];
                
                r_data[29621] <= r_data[29620];
                
                r_data[29622] <= r_data[29621];
                
                r_data[29623] <= r_data[29622];
                
                r_data[29624] <= r_data[29623];
                
                r_data[29625] <= r_data[29624];
                
                r_data[29626] <= r_data[29625];
                
                r_data[29627] <= r_data[29626];
                
                r_data[29628] <= r_data[29627];
                
                r_data[29629] <= r_data[29628];
                
                r_data[29630] <= r_data[29629];
                
                r_data[29631] <= r_data[29630];
                
                r_data[29632] <= r_data[29631];
                
                r_data[29633] <= r_data[29632];
                
                r_data[29634] <= r_data[29633];
                
                r_data[29635] <= r_data[29634];
                
                r_data[29636] <= r_data[29635];
                
                r_data[29637] <= r_data[29636];
                
                r_data[29638] <= r_data[29637];
                
                r_data[29639] <= r_data[29638];
                
                r_data[29640] <= r_data[29639];
                
                r_data[29641] <= r_data[29640];
                
                r_data[29642] <= r_data[29641];
                
                r_data[29643] <= r_data[29642];
                
                r_data[29644] <= r_data[29643];
                
                r_data[29645] <= r_data[29644];
                
                r_data[29646] <= r_data[29645];
                
                r_data[29647] <= r_data[29646];
                
                r_data[29648] <= r_data[29647];
                
                r_data[29649] <= r_data[29648];
                
                r_data[29650] <= r_data[29649];
                
                r_data[29651] <= r_data[29650];
                
                r_data[29652] <= r_data[29651];
                
                r_data[29653] <= r_data[29652];
                
                r_data[29654] <= r_data[29653];
                
                r_data[29655] <= r_data[29654];
                
                r_data[29656] <= r_data[29655];
                
                r_data[29657] <= r_data[29656];
                
                r_data[29658] <= r_data[29657];
                
                r_data[29659] <= r_data[29658];
                
                r_data[29660] <= r_data[29659];
                
                r_data[29661] <= r_data[29660];
                
                r_data[29662] <= r_data[29661];
                
                r_data[29663] <= r_data[29662];
                
                r_data[29664] <= r_data[29663];
                
                r_data[29665] <= r_data[29664];
                
                r_data[29666] <= r_data[29665];
                
                r_data[29667] <= r_data[29666];
                
                r_data[29668] <= r_data[29667];
                
                r_data[29669] <= r_data[29668];
                
                r_data[29670] <= r_data[29669];
                
                r_data[29671] <= r_data[29670];
                
                r_data[29672] <= r_data[29671];
                
                r_data[29673] <= r_data[29672];
                
                r_data[29674] <= r_data[29673];
                
                r_data[29675] <= r_data[29674];
                
                r_data[29676] <= r_data[29675];
                
                r_data[29677] <= r_data[29676];
                
                r_data[29678] <= r_data[29677];
                
                r_data[29679] <= r_data[29678];
                
                r_data[29680] <= r_data[29679];
                
                r_data[29681] <= r_data[29680];
                
                r_data[29682] <= r_data[29681];
                
                r_data[29683] <= r_data[29682];
                
                r_data[29684] <= r_data[29683];
                
                r_data[29685] <= r_data[29684];
                
                r_data[29686] <= r_data[29685];
                
                r_data[29687] <= r_data[29686];
                
                r_data[29688] <= r_data[29687];
                
                r_data[29689] <= r_data[29688];
                
                r_data[29690] <= r_data[29689];
                
                r_data[29691] <= r_data[29690];
                
                r_data[29692] <= r_data[29691];
                
                r_data[29693] <= r_data[29692];
                
                r_data[29694] <= r_data[29693];
                
                r_data[29695] <= r_data[29694];
                
                r_data[29696] <= r_data[29695];
                
                r_data[29697] <= r_data[29696];
                
                r_data[29698] <= r_data[29697];
                
                r_data[29699] <= r_data[29698];
                
                r_data[29700] <= r_data[29699];
                
                r_data[29701] <= r_data[29700];
                
                r_data[29702] <= r_data[29701];
                
                r_data[29703] <= r_data[29702];
                
                r_data[29704] <= r_data[29703];
                
                r_data[29705] <= r_data[29704];
                
                r_data[29706] <= r_data[29705];
                
                r_data[29707] <= r_data[29706];
                
                r_data[29708] <= r_data[29707];
                
                r_data[29709] <= r_data[29708];
                
                r_data[29710] <= r_data[29709];
                
                r_data[29711] <= r_data[29710];
                
                r_data[29712] <= r_data[29711];
                
                r_data[29713] <= r_data[29712];
                
                r_data[29714] <= r_data[29713];
                
                r_data[29715] <= r_data[29714];
                
                r_data[29716] <= r_data[29715];
                
                r_data[29717] <= r_data[29716];
                
                r_data[29718] <= r_data[29717];
                
                r_data[29719] <= r_data[29718];
                
                r_data[29720] <= r_data[29719];
                
                r_data[29721] <= r_data[29720];
                
                r_data[29722] <= r_data[29721];
                
                r_data[29723] <= r_data[29722];
                
                r_data[29724] <= r_data[29723];
                
                r_data[29725] <= r_data[29724];
                
                r_data[29726] <= r_data[29725];
                
                r_data[29727] <= r_data[29726];
                
                r_data[29728] <= r_data[29727];
                
                r_data[29729] <= r_data[29728];
                
                r_data[29730] <= r_data[29729];
                
                r_data[29731] <= r_data[29730];
                
                r_data[29732] <= r_data[29731];
                
                r_data[29733] <= r_data[29732];
                
                r_data[29734] <= r_data[29733];
                
                r_data[29735] <= r_data[29734];
                
                r_data[29736] <= r_data[29735];
                
                r_data[29737] <= r_data[29736];
                
                r_data[29738] <= r_data[29737];
                
                r_data[29739] <= r_data[29738];
                
                r_data[29740] <= r_data[29739];
                
                r_data[29741] <= r_data[29740];
                
                r_data[29742] <= r_data[29741];
                
                r_data[29743] <= r_data[29742];
                
                r_data[29744] <= r_data[29743];
                
                r_data[29745] <= r_data[29744];
                
                r_data[29746] <= r_data[29745];
                
                r_data[29747] <= r_data[29746];
                
                r_data[29748] <= r_data[29747];
                
                r_data[29749] <= r_data[29748];
                
                r_data[29750] <= r_data[29749];
                
                r_data[29751] <= r_data[29750];
                
                r_data[29752] <= r_data[29751];
                
                r_data[29753] <= r_data[29752];
                
                r_data[29754] <= r_data[29753];
                
                r_data[29755] <= r_data[29754];
                
                r_data[29756] <= r_data[29755];
                
                r_data[29757] <= r_data[29756];
                
                r_data[29758] <= r_data[29757];
                
                r_data[29759] <= r_data[29758];
                
                r_data[29760] <= r_data[29759];
                
                r_data[29761] <= r_data[29760];
                
                r_data[29762] <= r_data[29761];
                
                r_data[29763] <= r_data[29762];
                
                r_data[29764] <= r_data[29763];
                
                r_data[29765] <= r_data[29764];
                
                r_data[29766] <= r_data[29765];
                
                r_data[29767] <= r_data[29766];
                
                r_data[29768] <= r_data[29767];
                
                r_data[29769] <= r_data[29768];
                
                r_data[29770] <= r_data[29769];
                
                r_data[29771] <= r_data[29770];
                
                r_data[29772] <= r_data[29771];
                
                r_data[29773] <= r_data[29772];
                
                r_data[29774] <= r_data[29773];
                
                r_data[29775] <= r_data[29774];
                
                r_data[29776] <= r_data[29775];
                
                r_data[29777] <= r_data[29776];
                
                r_data[29778] <= r_data[29777];
                
                r_data[29779] <= r_data[29778];
                
                r_data[29780] <= r_data[29779];
                
                r_data[29781] <= r_data[29780];
                
                r_data[29782] <= r_data[29781];
                
                r_data[29783] <= r_data[29782];
                
                r_data[29784] <= r_data[29783];
                
                r_data[29785] <= r_data[29784];
                
                r_data[29786] <= r_data[29785];
                
                r_data[29787] <= r_data[29786];
                
                r_data[29788] <= r_data[29787];
                
                r_data[29789] <= r_data[29788];
                
                r_data[29790] <= r_data[29789];
                
                r_data[29791] <= r_data[29790];
                
                r_data[29792] <= r_data[29791];
                
                r_data[29793] <= r_data[29792];
                
                r_data[29794] <= r_data[29793];
                
                r_data[29795] <= r_data[29794];
                
                r_data[29796] <= r_data[29795];
                
                r_data[29797] <= r_data[29796];
                
                r_data[29798] <= r_data[29797];
                
                r_data[29799] <= r_data[29798];
                
                r_data[29800] <= r_data[29799];
                
                r_data[29801] <= r_data[29800];
                
                r_data[29802] <= r_data[29801];
                
                r_data[29803] <= r_data[29802];
                
                r_data[29804] <= r_data[29803];
                
                r_data[29805] <= r_data[29804];
                
                r_data[29806] <= r_data[29805];
                
                r_data[29807] <= r_data[29806];
                
                r_data[29808] <= r_data[29807];
                
                r_data[29809] <= r_data[29808];
                
                r_data[29810] <= r_data[29809];
                
                r_data[29811] <= r_data[29810];
                
                r_data[29812] <= r_data[29811];
                
                r_data[29813] <= r_data[29812];
                
                r_data[29814] <= r_data[29813];
                
                r_data[29815] <= r_data[29814];
                
                r_data[29816] <= r_data[29815];
                
                r_data[29817] <= r_data[29816];
                
                r_data[29818] <= r_data[29817];
                
                r_data[29819] <= r_data[29818];
                
                r_data[29820] <= r_data[29819];
                
                r_data[29821] <= r_data[29820];
                
                r_data[29822] <= r_data[29821];
                
                r_data[29823] <= r_data[29822];
                
                r_data[29824] <= r_data[29823];
                
                r_data[29825] <= r_data[29824];
                
                r_data[29826] <= r_data[29825];
                
                r_data[29827] <= r_data[29826];
                
                r_data[29828] <= r_data[29827];
                
                r_data[29829] <= r_data[29828];
                
                r_data[29830] <= r_data[29829];
                
                r_data[29831] <= r_data[29830];
                
                r_data[29832] <= r_data[29831];
                
                r_data[29833] <= r_data[29832];
                
                r_data[29834] <= r_data[29833];
                
                r_data[29835] <= r_data[29834];
                
                r_data[29836] <= r_data[29835];
                
                r_data[29837] <= r_data[29836];
                
                r_data[29838] <= r_data[29837];
                
                r_data[29839] <= r_data[29838];
                
                r_data[29840] <= r_data[29839];
                
                r_data[29841] <= r_data[29840];
                
                r_data[29842] <= r_data[29841];
                
                r_data[29843] <= r_data[29842];
                
                r_data[29844] <= r_data[29843];
                
                r_data[29845] <= r_data[29844];
                
                r_data[29846] <= r_data[29845];
                
                r_data[29847] <= r_data[29846];
                
                r_data[29848] <= r_data[29847];
                
                r_data[29849] <= r_data[29848];
                
                r_data[29850] <= r_data[29849];
                
                r_data[29851] <= r_data[29850];
                
                r_data[29852] <= r_data[29851];
                
                r_data[29853] <= r_data[29852];
                
                r_data[29854] <= r_data[29853];
                
                r_data[29855] <= r_data[29854];
                
                r_data[29856] <= r_data[29855];
                
                r_data[29857] <= r_data[29856];
                
                r_data[29858] <= r_data[29857];
                
                r_data[29859] <= r_data[29858];
                
                r_data[29860] <= r_data[29859];
                
                r_data[29861] <= r_data[29860];
                
                r_data[29862] <= r_data[29861];
                
                r_data[29863] <= r_data[29862];
                
                r_data[29864] <= r_data[29863];
                
                r_data[29865] <= r_data[29864];
                
                r_data[29866] <= r_data[29865];
                
                r_data[29867] <= r_data[29866];
                
                r_data[29868] <= r_data[29867];
                
                r_data[29869] <= r_data[29868];
                
                r_data[29870] <= r_data[29869];
                
                r_data[29871] <= r_data[29870];
                
                r_data[29872] <= r_data[29871];
                
                r_data[29873] <= r_data[29872];
                
                r_data[29874] <= r_data[29873];
                
                r_data[29875] <= r_data[29874];
                
                r_data[29876] <= r_data[29875];
                
                r_data[29877] <= r_data[29876];
                
                r_data[29878] <= r_data[29877];
                
                r_data[29879] <= r_data[29878];
                
                r_data[29880] <= r_data[29879];
                
                r_data[29881] <= r_data[29880];
                
                r_data[29882] <= r_data[29881];
                
                r_data[29883] <= r_data[29882];
                
                r_data[29884] <= r_data[29883];
                
                r_data[29885] <= r_data[29884];
                
                r_data[29886] <= r_data[29885];
                
                r_data[29887] <= r_data[29886];
                
                r_data[29888] <= r_data[29887];
                
                r_data[29889] <= r_data[29888];
                
                r_data[29890] <= r_data[29889];
                
                r_data[29891] <= r_data[29890];
                
                r_data[29892] <= r_data[29891];
                
                r_data[29893] <= r_data[29892];
                
                r_data[29894] <= r_data[29893];
                
                r_data[29895] <= r_data[29894];
                
                r_data[29896] <= r_data[29895];
                
                r_data[29897] <= r_data[29896];
                
                r_data[29898] <= r_data[29897];
                
                r_data[29899] <= r_data[29898];
                
                r_data[29900] <= r_data[29899];
                
                r_data[29901] <= r_data[29900];
                
                r_data[29902] <= r_data[29901];
                
                r_data[29903] <= r_data[29902];
                
                r_data[29904] <= r_data[29903];
                
                r_data[29905] <= r_data[29904];
                
                r_data[29906] <= r_data[29905];
                
                r_data[29907] <= r_data[29906];
                
                r_data[29908] <= r_data[29907];
                
                r_data[29909] <= r_data[29908];
                
                r_data[29910] <= r_data[29909];
                
                r_data[29911] <= r_data[29910];
                
                r_data[29912] <= r_data[29911];
                
                r_data[29913] <= r_data[29912];
                
                r_data[29914] <= r_data[29913];
                
                r_data[29915] <= r_data[29914];
                
                r_data[29916] <= r_data[29915];
                
                r_data[29917] <= r_data[29916];
                
                r_data[29918] <= r_data[29917];
                
                r_data[29919] <= r_data[29918];
                
                r_data[29920] <= r_data[29919];
                
                r_data[29921] <= r_data[29920];
                
                r_data[29922] <= r_data[29921];
                
                r_data[29923] <= r_data[29922];
                
                r_data[29924] <= r_data[29923];
                
                r_data[29925] <= r_data[29924];
                
                r_data[29926] <= r_data[29925];
                
                r_data[29927] <= r_data[29926];
                
                r_data[29928] <= r_data[29927];
                
                r_data[29929] <= r_data[29928];
                
                r_data[29930] <= r_data[29929];
                
                r_data[29931] <= r_data[29930];
                
                r_data[29932] <= r_data[29931];
                
                r_data[29933] <= r_data[29932];
                
                r_data[29934] <= r_data[29933];
                
                r_data[29935] <= r_data[29934];
                
                r_data[29936] <= r_data[29935];
                
                r_data[29937] <= r_data[29936];
                
                r_data[29938] <= r_data[29937];
                
                r_data[29939] <= r_data[29938];
                
                r_data[29940] <= r_data[29939];
                
                r_data[29941] <= r_data[29940];
                
                r_data[29942] <= r_data[29941];
                
                r_data[29943] <= r_data[29942];
                
                r_data[29944] <= r_data[29943];
                
                r_data[29945] <= r_data[29944];
                
                r_data[29946] <= r_data[29945];
                
                r_data[29947] <= r_data[29946];
                
                r_data[29948] <= r_data[29947];
                
                r_data[29949] <= r_data[29948];
                
                r_data[29950] <= r_data[29949];
                
                r_data[29951] <= r_data[29950];
                
                r_data[29952] <= r_data[29951];
                
                r_data[29953] <= r_data[29952];
                
                r_data[29954] <= r_data[29953];
                
                r_data[29955] <= r_data[29954];
                
                r_data[29956] <= r_data[29955];
                
                r_data[29957] <= r_data[29956];
                
                r_data[29958] <= r_data[29957];
                
                r_data[29959] <= r_data[29958];
                
                r_data[29960] <= r_data[29959];
                
                r_data[29961] <= r_data[29960];
                
                r_data[29962] <= r_data[29961];
                
                r_data[29963] <= r_data[29962];
                
                r_data[29964] <= r_data[29963];
                
                r_data[29965] <= r_data[29964];
                
                r_data[29966] <= r_data[29965];
                
                r_data[29967] <= r_data[29966];
                
                r_data[29968] <= r_data[29967];
                
                r_data[29969] <= r_data[29968];
                
                r_data[29970] <= r_data[29969];
                
                r_data[29971] <= r_data[29970];
                
                r_data[29972] <= r_data[29971];
                
                r_data[29973] <= r_data[29972];
                
                r_data[29974] <= r_data[29973];
                
                r_data[29975] <= r_data[29974];
                
                r_data[29976] <= r_data[29975];
                
                r_data[29977] <= r_data[29976];
                
                r_data[29978] <= r_data[29977];
                
                r_data[29979] <= r_data[29978];
                
                r_data[29980] <= r_data[29979];
                
                r_data[29981] <= r_data[29980];
                
                r_data[29982] <= r_data[29981];
                
                r_data[29983] <= r_data[29982];
                
                r_data[29984] <= r_data[29983];
                
                r_data[29985] <= r_data[29984];
                
                r_data[29986] <= r_data[29985];
                
                r_data[29987] <= r_data[29986];
                
                r_data[29988] <= r_data[29987];
                
                r_data[29989] <= r_data[29988];
                
                r_data[29990] <= r_data[29989];
                
                r_data[29991] <= r_data[29990];
                
                r_data[29992] <= r_data[29991];
                
                r_data[29993] <= r_data[29992];
                
                r_data[29994] <= r_data[29993];
                
                r_data[29995] <= r_data[29994];
                
                r_data[29996] <= r_data[29995];
                
                r_data[29997] <= r_data[29996];
                
                r_data[29998] <= r_data[29997];
                
                r_data[29999] <= r_data[29998];
                
                r_data[30000] <= r_data[29999];
                
                r_data[30001] <= r_data[30000];
                
                r_data[30002] <= r_data[30001];
                
                r_data[30003] <= r_data[30002];
                
                r_data[30004] <= r_data[30003];
                
                r_data[30005] <= r_data[30004];
                
                r_data[30006] <= r_data[30005];
                
                r_data[30007] <= r_data[30006];
                
                r_data[30008] <= r_data[30007];
                
                r_data[30009] <= r_data[30008];
                
                r_data[30010] <= r_data[30009];
                
                r_data[30011] <= r_data[30010];
                
                r_data[30012] <= r_data[30011];
                
                r_data[30013] <= r_data[30012];
                
                r_data[30014] <= r_data[30013];
                
                r_data[30015] <= r_data[30014];
                
                r_data[30016] <= r_data[30015];
                
                r_data[30017] <= r_data[30016];
                
                r_data[30018] <= r_data[30017];
                
                r_data[30019] <= r_data[30018];
                
                r_data[30020] <= r_data[30019];
                
                r_data[30021] <= r_data[30020];
                
                r_data[30022] <= r_data[30021];
                
                r_data[30023] <= r_data[30022];
                
                r_data[30024] <= r_data[30023];
                
                r_data[30025] <= r_data[30024];
                
                r_data[30026] <= r_data[30025];
                
                r_data[30027] <= r_data[30026];
                
                r_data[30028] <= r_data[30027];
                
                r_data[30029] <= r_data[30028];
                
                r_data[30030] <= r_data[30029];
                
                r_data[30031] <= r_data[30030];
                
                r_data[30032] <= r_data[30031];
                
                r_data[30033] <= r_data[30032];
                
                r_data[30034] <= r_data[30033];
                
                r_data[30035] <= r_data[30034];
                
                r_data[30036] <= r_data[30035];
                
                r_data[30037] <= r_data[30036];
                
                r_data[30038] <= r_data[30037];
                
                r_data[30039] <= r_data[30038];
                
                r_data[30040] <= r_data[30039];
                
                r_data[30041] <= r_data[30040];
                
                r_data[30042] <= r_data[30041];
                
                r_data[30043] <= r_data[30042];
                
                r_data[30044] <= r_data[30043];
                
                r_data[30045] <= r_data[30044];
                
                r_data[30046] <= r_data[30045];
                
                r_data[30047] <= r_data[30046];
                
                r_data[30048] <= r_data[30047];
                
                r_data[30049] <= r_data[30048];
                
                r_data[30050] <= r_data[30049];
                
                r_data[30051] <= r_data[30050];
                
                r_data[30052] <= r_data[30051];
                
                r_data[30053] <= r_data[30052];
                
                r_data[30054] <= r_data[30053];
                
                r_data[30055] <= r_data[30054];
                
                r_data[30056] <= r_data[30055];
                
                r_data[30057] <= r_data[30056];
                
                r_data[30058] <= r_data[30057];
                
                r_data[30059] <= r_data[30058];
                
                r_data[30060] <= r_data[30059];
                
                r_data[30061] <= r_data[30060];
                
                r_data[30062] <= r_data[30061];
                
                r_data[30063] <= r_data[30062];
                
                r_data[30064] <= r_data[30063];
                
                r_data[30065] <= r_data[30064];
                
                r_data[30066] <= r_data[30065];
                
                r_data[30067] <= r_data[30066];
                
                r_data[30068] <= r_data[30067];
                
                r_data[30069] <= r_data[30068];
                
                r_data[30070] <= r_data[30069];
                
                r_data[30071] <= r_data[30070];
                
                r_data[30072] <= r_data[30071];
                
                r_data[30073] <= r_data[30072];
                
                r_data[30074] <= r_data[30073];
                
                r_data[30075] <= r_data[30074];
                
                r_data[30076] <= r_data[30075];
                
                r_data[30077] <= r_data[30076];
                
                r_data[30078] <= r_data[30077];
                
                r_data[30079] <= r_data[30078];
                
                r_data[30080] <= r_data[30079];
                
                r_data[30081] <= r_data[30080];
                
                r_data[30082] <= r_data[30081];
                
                r_data[30083] <= r_data[30082];
                
                r_data[30084] <= r_data[30083];
                
                r_data[30085] <= r_data[30084];
                
                r_data[30086] <= r_data[30085];
                
                r_data[30087] <= r_data[30086];
                
                r_data[30088] <= r_data[30087];
                
                r_data[30089] <= r_data[30088];
                
                r_data[30090] <= r_data[30089];
                
                r_data[30091] <= r_data[30090];
                
                r_data[30092] <= r_data[30091];
                
                r_data[30093] <= r_data[30092];
                
                r_data[30094] <= r_data[30093];
                
                r_data[30095] <= r_data[30094];
                
                r_data[30096] <= r_data[30095];
                
                r_data[30097] <= r_data[30096];
                
                r_data[30098] <= r_data[30097];
                
                r_data[30099] <= r_data[30098];
                
                r_data[30100] <= r_data[30099];
                
                r_data[30101] <= r_data[30100];
                
                r_data[30102] <= r_data[30101];
                
                r_data[30103] <= r_data[30102];
                
                r_data[30104] <= r_data[30103];
                
                r_data[30105] <= r_data[30104];
                
                r_data[30106] <= r_data[30105];
                
                r_data[30107] <= r_data[30106];
                
                r_data[30108] <= r_data[30107];
                
                r_data[30109] <= r_data[30108];
                
                r_data[30110] <= r_data[30109];
                
                r_data[30111] <= r_data[30110];
                
                r_data[30112] <= r_data[30111];
                
                r_data[30113] <= r_data[30112];
                
                r_data[30114] <= r_data[30113];
                
                r_data[30115] <= r_data[30114];
                
                r_data[30116] <= r_data[30115];
                
                r_data[30117] <= r_data[30116];
                
                r_data[30118] <= r_data[30117];
                
                r_data[30119] <= r_data[30118];
                
                r_data[30120] <= r_data[30119];
                
                r_data[30121] <= r_data[30120];
                
                r_data[30122] <= r_data[30121];
                
                r_data[30123] <= r_data[30122];
                
                r_data[30124] <= r_data[30123];
                
                r_data[30125] <= r_data[30124];
                
                r_data[30126] <= r_data[30125];
                
                r_data[30127] <= r_data[30126];
                
                r_data[30128] <= r_data[30127];
                
                r_data[30129] <= r_data[30128];
                
                r_data[30130] <= r_data[30129];
                
                r_data[30131] <= r_data[30130];
                
                r_data[30132] <= r_data[30131];
                
                r_data[30133] <= r_data[30132];
                
                r_data[30134] <= r_data[30133];
                
                r_data[30135] <= r_data[30134];
                
                r_data[30136] <= r_data[30135];
                
                r_data[30137] <= r_data[30136];
                
                r_data[30138] <= r_data[30137];
                
                r_data[30139] <= r_data[30138];
                
                r_data[30140] <= r_data[30139];
                
                r_data[30141] <= r_data[30140];
                
                r_data[30142] <= r_data[30141];
                
                r_data[30143] <= r_data[30142];
                
                r_data[30144] <= r_data[30143];
                
                r_data[30145] <= r_data[30144];
                
                r_data[30146] <= r_data[30145];
                
                r_data[30147] <= r_data[30146];
                
                r_data[30148] <= r_data[30147];
                
                r_data[30149] <= r_data[30148];
                
                r_data[30150] <= r_data[30149];
                
                r_data[30151] <= r_data[30150];
                
                r_data[30152] <= r_data[30151];
                
                r_data[30153] <= r_data[30152];
                
                r_data[30154] <= r_data[30153];
                
                r_data[30155] <= r_data[30154];
                
                r_data[30156] <= r_data[30155];
                
                r_data[30157] <= r_data[30156];
                
                r_data[30158] <= r_data[30157];
                
                r_data[30159] <= r_data[30158];
                
                r_data[30160] <= r_data[30159];
                
                r_data[30161] <= r_data[30160];
                
                r_data[30162] <= r_data[30161];
                
                r_data[30163] <= r_data[30162];
                
                r_data[30164] <= r_data[30163];
                
                r_data[30165] <= r_data[30164];
                
                r_data[30166] <= r_data[30165];
                
                r_data[30167] <= r_data[30166];
                
                r_data[30168] <= r_data[30167];
                
                r_data[30169] <= r_data[30168];
                
                r_data[30170] <= r_data[30169];
                
                r_data[30171] <= r_data[30170];
                
                r_data[30172] <= r_data[30171];
                
                r_data[30173] <= r_data[30172];
                
                r_data[30174] <= r_data[30173];
                
                r_data[30175] <= r_data[30174];
                
                r_data[30176] <= r_data[30175];
                
                r_data[30177] <= r_data[30176];
                
                r_data[30178] <= r_data[30177];
                
                r_data[30179] <= r_data[30178];
                
                r_data[30180] <= r_data[30179];
                
                r_data[30181] <= r_data[30180];
                
                r_data[30182] <= r_data[30181];
                
                r_data[30183] <= r_data[30182];
                
                r_data[30184] <= r_data[30183];
                
                r_data[30185] <= r_data[30184];
                
                r_data[30186] <= r_data[30185];
                
                r_data[30187] <= r_data[30186];
                
                r_data[30188] <= r_data[30187];
                
                r_data[30189] <= r_data[30188];
                
                r_data[30190] <= r_data[30189];
                
                r_data[30191] <= r_data[30190];
                
                r_data[30192] <= r_data[30191];
                
                r_data[30193] <= r_data[30192];
                
                r_data[30194] <= r_data[30193];
                
                r_data[30195] <= r_data[30194];
                
                r_data[30196] <= r_data[30195];
                
                r_data[30197] <= r_data[30196];
                
                r_data[30198] <= r_data[30197];
                
                r_data[30199] <= r_data[30198];
                
                r_data[30200] <= r_data[30199];
                
                r_data[30201] <= r_data[30200];
                
                r_data[30202] <= r_data[30201];
                
                r_data[30203] <= r_data[30202];
                
                r_data[30204] <= r_data[30203];
                
                r_data[30205] <= r_data[30204];
                
                r_data[30206] <= r_data[30205];
                
                r_data[30207] <= r_data[30206];
                
                r_data[30208] <= r_data[30207];
                
                r_data[30209] <= r_data[30208];
                
                r_data[30210] <= r_data[30209];
                
                r_data[30211] <= r_data[30210];
                
                r_data[30212] <= r_data[30211];
                
                r_data[30213] <= r_data[30212];
                
                r_data[30214] <= r_data[30213];
                
                r_data[30215] <= r_data[30214];
                
                r_data[30216] <= r_data[30215];
                
                r_data[30217] <= r_data[30216];
                
                r_data[30218] <= r_data[30217];
                
                r_data[30219] <= r_data[30218];
                
                r_data[30220] <= r_data[30219];
                
                r_data[30221] <= r_data[30220];
                
                r_data[30222] <= r_data[30221];
                
                r_data[30223] <= r_data[30222];
                
                r_data[30224] <= r_data[30223];
                
                r_data[30225] <= r_data[30224];
                
                r_data[30226] <= r_data[30225];
                
                r_data[30227] <= r_data[30226];
                
                r_data[30228] <= r_data[30227];
                
                r_data[30229] <= r_data[30228];
                
                r_data[30230] <= r_data[30229];
                
                r_data[30231] <= r_data[30230];
                
                r_data[30232] <= r_data[30231];
                
                r_data[30233] <= r_data[30232];
                
                r_data[30234] <= r_data[30233];
                
                r_data[30235] <= r_data[30234];
                
                r_data[30236] <= r_data[30235];
                
                r_data[30237] <= r_data[30236];
                
                r_data[30238] <= r_data[30237];
                
                r_data[30239] <= r_data[30238];
                
                r_data[30240] <= r_data[30239];
                
                r_data[30241] <= r_data[30240];
                
                r_data[30242] <= r_data[30241];
                
                r_data[30243] <= r_data[30242];
                
                r_data[30244] <= r_data[30243];
                
                r_data[30245] <= r_data[30244];
                
                r_data[30246] <= r_data[30245];
                
                r_data[30247] <= r_data[30246];
                
                r_data[30248] <= r_data[30247];
                
                r_data[30249] <= r_data[30248];
                
                r_data[30250] <= r_data[30249];
                
                r_data[30251] <= r_data[30250];
                
                r_data[30252] <= r_data[30251];
                
                r_data[30253] <= r_data[30252];
                
                r_data[30254] <= r_data[30253];
                
                r_data[30255] <= r_data[30254];
                
                r_data[30256] <= r_data[30255];
                
                r_data[30257] <= r_data[30256];
                
                r_data[30258] <= r_data[30257];
                
                r_data[30259] <= r_data[30258];
                
                r_data[30260] <= r_data[30259];
                
                r_data[30261] <= r_data[30260];
                
                r_data[30262] <= r_data[30261];
                
                r_data[30263] <= r_data[30262];
                
                r_data[30264] <= r_data[30263];
                
                r_data[30265] <= r_data[30264];
                
                r_data[30266] <= r_data[30265];
                
                r_data[30267] <= r_data[30266];
                
                r_data[30268] <= r_data[30267];
                
                r_data[30269] <= r_data[30268];
                
                r_data[30270] <= r_data[30269];
                
                r_data[30271] <= r_data[30270];
                
                r_data[30272] <= r_data[30271];
                
                r_data[30273] <= r_data[30272];
                
                r_data[30274] <= r_data[30273];
                
                r_data[30275] <= r_data[30274];
                
                r_data[30276] <= r_data[30275];
                
                r_data[30277] <= r_data[30276];
                
                r_data[30278] <= r_data[30277];
                
                r_data[30279] <= r_data[30278];
                
                r_data[30280] <= r_data[30279];
                
                r_data[30281] <= r_data[30280];
                
                r_data[30282] <= r_data[30281];
                
                r_data[30283] <= r_data[30282];
                
                r_data[30284] <= r_data[30283];
                
                r_data[30285] <= r_data[30284];
                
                r_data[30286] <= r_data[30285];
                
                r_data[30287] <= r_data[30286];
                
                r_data[30288] <= r_data[30287];
                
                r_data[30289] <= r_data[30288];
                
                r_data[30290] <= r_data[30289];
                
                r_data[30291] <= r_data[30290];
                
                r_data[30292] <= r_data[30291];
                
                r_data[30293] <= r_data[30292];
                
                r_data[30294] <= r_data[30293];
                
                r_data[30295] <= r_data[30294];
                
                r_data[30296] <= r_data[30295];
                
                r_data[30297] <= r_data[30296];
                
                r_data[30298] <= r_data[30297];
                
                r_data[30299] <= r_data[30298];
                
                r_data[30300] <= r_data[30299];
                
                r_data[30301] <= r_data[30300];
                
                r_data[30302] <= r_data[30301];
                
                r_data[30303] <= r_data[30302];
                
                r_data[30304] <= r_data[30303];
                
                r_data[30305] <= r_data[30304];
                
                r_data[30306] <= r_data[30305];
                
                r_data[30307] <= r_data[30306];
                
                r_data[30308] <= r_data[30307];
                
                r_data[30309] <= r_data[30308];
                
                r_data[30310] <= r_data[30309];
                
                r_data[30311] <= r_data[30310];
                
                r_data[30312] <= r_data[30311];
                
                r_data[30313] <= r_data[30312];
                
                r_data[30314] <= r_data[30313];
                
                r_data[30315] <= r_data[30314];
                
                r_data[30316] <= r_data[30315];
                
                r_data[30317] <= r_data[30316];
                
                r_data[30318] <= r_data[30317];
                
                r_data[30319] <= r_data[30318];
                
                r_data[30320] <= r_data[30319];
                
                r_data[30321] <= r_data[30320];
                
                r_data[30322] <= r_data[30321];
                
                r_data[30323] <= r_data[30322];
                
                r_data[30324] <= r_data[30323];
                
                r_data[30325] <= r_data[30324];
                
                r_data[30326] <= r_data[30325];
                
                r_data[30327] <= r_data[30326];
                
                r_data[30328] <= r_data[30327];
                
                r_data[30329] <= r_data[30328];
                
                r_data[30330] <= r_data[30329];
                
                r_data[30331] <= r_data[30330];
                
                r_data[30332] <= r_data[30331];
                
                r_data[30333] <= r_data[30332];
                
                r_data[30334] <= r_data[30333];
                
                r_data[30335] <= r_data[30334];
                
                r_data[30336] <= r_data[30335];
                
                r_data[30337] <= r_data[30336];
                
                r_data[30338] <= r_data[30337];
                
                r_data[30339] <= r_data[30338];
                
                r_data[30340] <= r_data[30339];
                
                r_data[30341] <= r_data[30340];
                
                r_data[30342] <= r_data[30341];
                
                r_data[30343] <= r_data[30342];
                
                r_data[30344] <= r_data[30343];
                
                r_data[30345] <= r_data[30344];
                
                r_data[30346] <= r_data[30345];
                
                r_data[30347] <= r_data[30346];
                
                r_data[30348] <= r_data[30347];
                
                r_data[30349] <= r_data[30348];
                
                r_data[30350] <= r_data[30349];
                
                r_data[30351] <= r_data[30350];
                
                r_data[30352] <= r_data[30351];
                
                r_data[30353] <= r_data[30352];
                
                r_data[30354] <= r_data[30353];
                
                r_data[30355] <= r_data[30354];
                
                r_data[30356] <= r_data[30355];
                
                r_data[30357] <= r_data[30356];
                
                r_data[30358] <= r_data[30357];
                
                r_data[30359] <= r_data[30358];
                
                r_data[30360] <= r_data[30359];
                
                r_data[30361] <= r_data[30360];
                
                r_data[30362] <= r_data[30361];
                
                r_data[30363] <= r_data[30362];
                
                r_data[30364] <= r_data[30363];
                
                r_data[30365] <= r_data[30364];
                
                r_data[30366] <= r_data[30365];
                
                r_data[30367] <= r_data[30366];
                
                r_data[30368] <= r_data[30367];
                
                r_data[30369] <= r_data[30368];
                
                r_data[30370] <= r_data[30369];
                
                r_data[30371] <= r_data[30370];
                
                r_data[30372] <= r_data[30371];
                
                r_data[30373] <= r_data[30372];
                
                r_data[30374] <= r_data[30373];
                
                r_data[30375] <= r_data[30374];
                
                r_data[30376] <= r_data[30375];
                
                r_data[30377] <= r_data[30376];
                
                r_data[30378] <= r_data[30377];
                
                r_data[30379] <= r_data[30378];
                
                r_data[30380] <= r_data[30379];
                
                r_data[30381] <= r_data[30380];
                
                r_data[30382] <= r_data[30381];
                
                r_data[30383] <= r_data[30382];
                
                r_data[30384] <= r_data[30383];
                
                r_data[30385] <= r_data[30384];
                
                r_data[30386] <= r_data[30385];
                
                r_data[30387] <= r_data[30386];
                
                r_data[30388] <= r_data[30387];
                
                r_data[30389] <= r_data[30388];
                
                r_data[30390] <= r_data[30389];
                
                r_data[30391] <= r_data[30390];
                
                r_data[30392] <= r_data[30391];
                
                r_data[30393] <= r_data[30392];
                
                r_data[30394] <= r_data[30393];
                
                r_data[30395] <= r_data[30394];
                
                r_data[30396] <= r_data[30395];
                
                r_data[30397] <= r_data[30396];
                
                r_data[30398] <= r_data[30397];
                
                r_data[30399] <= r_data[30398];
                
                r_data[30400] <= r_data[30399];
                
                r_data[30401] <= r_data[30400];
                
                r_data[30402] <= r_data[30401];
                
                r_data[30403] <= r_data[30402];
                
                r_data[30404] <= r_data[30403];
                
                r_data[30405] <= r_data[30404];
                
                r_data[30406] <= r_data[30405];
                
                r_data[30407] <= r_data[30406];
                
                r_data[30408] <= r_data[30407];
                
                r_data[30409] <= r_data[30408];
                
                r_data[30410] <= r_data[30409];
                
                r_data[30411] <= r_data[30410];
                
                r_data[30412] <= r_data[30411];
                
                r_data[30413] <= r_data[30412];
                
                r_data[30414] <= r_data[30413];
                
                r_data[30415] <= r_data[30414];
                
                r_data[30416] <= r_data[30415];
                
                r_data[30417] <= r_data[30416];
                
                r_data[30418] <= r_data[30417];
                
                r_data[30419] <= r_data[30418];
                
                r_data[30420] <= r_data[30419];
                
                r_data[30421] <= r_data[30420];
                
                r_data[30422] <= r_data[30421];
                
                r_data[30423] <= r_data[30422];
                
                r_data[30424] <= r_data[30423];
                
                r_data[30425] <= r_data[30424];
                
                r_data[30426] <= r_data[30425];
                
                r_data[30427] <= r_data[30426];
                
                r_data[30428] <= r_data[30427];
                
                r_data[30429] <= r_data[30428];
                
                r_data[30430] <= r_data[30429];
                
                r_data[30431] <= r_data[30430];
                
                r_data[30432] <= r_data[30431];
                
                r_data[30433] <= r_data[30432];
                
                r_data[30434] <= r_data[30433];
                
                r_data[30435] <= r_data[30434];
                
                r_data[30436] <= r_data[30435];
                
                r_data[30437] <= r_data[30436];
                
                r_data[30438] <= r_data[30437];
                
                r_data[30439] <= r_data[30438];
                
                r_data[30440] <= r_data[30439];
                
                r_data[30441] <= r_data[30440];
                
                r_data[30442] <= r_data[30441];
                
                r_data[30443] <= r_data[30442];
                
                r_data[30444] <= r_data[30443];
                
                r_data[30445] <= r_data[30444];
                
                r_data[30446] <= r_data[30445];
                
                r_data[30447] <= r_data[30446];
                
                r_data[30448] <= r_data[30447];
                
                r_data[30449] <= r_data[30448];
                
                r_data[30450] <= r_data[30449];
                
                r_data[30451] <= r_data[30450];
                
                r_data[30452] <= r_data[30451];
                
                r_data[30453] <= r_data[30452];
                
                r_data[30454] <= r_data[30453];
                
                r_data[30455] <= r_data[30454];
                
                r_data[30456] <= r_data[30455];
                
                r_data[30457] <= r_data[30456];
                
                r_data[30458] <= r_data[30457];
                
                r_data[30459] <= r_data[30458];
                
                r_data[30460] <= r_data[30459];
                
                r_data[30461] <= r_data[30460];
                
                r_data[30462] <= r_data[30461];
                
                r_data[30463] <= r_data[30462];
                
                r_data[30464] <= r_data[30463];
                
                r_data[30465] <= r_data[30464];
                
                r_data[30466] <= r_data[30465];
                
                r_data[30467] <= r_data[30466];
                
                r_data[30468] <= r_data[30467];
                
                r_data[30469] <= r_data[30468];
                
                r_data[30470] <= r_data[30469];
                
                r_data[30471] <= r_data[30470];
                
                r_data[30472] <= r_data[30471];
                
                r_data[30473] <= r_data[30472];
                
                r_data[30474] <= r_data[30473];
                
                r_data[30475] <= r_data[30474];
                
                r_data[30476] <= r_data[30475];
                
                r_data[30477] <= r_data[30476];
                
                r_data[30478] <= r_data[30477];
                
                r_data[30479] <= r_data[30478];
                
                r_data[30480] <= r_data[30479];
                
                r_data[30481] <= r_data[30480];
                
                r_data[30482] <= r_data[30481];
                
                r_data[30483] <= r_data[30482];
                
                r_data[30484] <= r_data[30483];
                
                r_data[30485] <= r_data[30484];
                
                r_data[30486] <= r_data[30485];
                
                r_data[30487] <= r_data[30486];
                
                r_data[30488] <= r_data[30487];
                
                r_data[30489] <= r_data[30488];
                
                r_data[30490] <= r_data[30489];
                
                r_data[30491] <= r_data[30490];
                
                r_data[30492] <= r_data[30491];
                
                r_data[30493] <= r_data[30492];
                
                r_data[30494] <= r_data[30493];
                
                r_data[30495] <= r_data[30494];
                
                r_data[30496] <= r_data[30495];
                
                r_data[30497] <= r_data[30496];
                
                r_data[30498] <= r_data[30497];
                
                r_data[30499] <= r_data[30498];
                
                r_data[30500] <= r_data[30499];
                
                r_data[30501] <= r_data[30500];
                
                r_data[30502] <= r_data[30501];
                
                r_data[30503] <= r_data[30502];
                
                r_data[30504] <= r_data[30503];
                
                r_data[30505] <= r_data[30504];
                
                r_data[30506] <= r_data[30505];
                
                r_data[30507] <= r_data[30506];
                
                r_data[30508] <= r_data[30507];
                
                r_data[30509] <= r_data[30508];
                
                r_data[30510] <= r_data[30509];
                
                r_data[30511] <= r_data[30510];
                
                r_data[30512] <= r_data[30511];
                
                r_data[30513] <= r_data[30512];
                
                r_data[30514] <= r_data[30513];
                
                r_data[30515] <= r_data[30514];
                
                r_data[30516] <= r_data[30515];
                
                r_data[30517] <= r_data[30516];
                
                r_data[30518] <= r_data[30517];
                
                r_data[30519] <= r_data[30518];
                
                r_data[30520] <= r_data[30519];
                
                r_data[30521] <= r_data[30520];
                
                r_data[30522] <= r_data[30521];
                
                r_data[30523] <= r_data[30522];
                
                r_data[30524] <= r_data[30523];
                
                r_data[30525] <= r_data[30524];
                
                r_data[30526] <= r_data[30525];
                
                r_data[30527] <= r_data[30526];
                
                r_data[30528] <= r_data[30527];
                
                r_data[30529] <= r_data[30528];
                
                r_data[30530] <= r_data[30529];
                
                r_data[30531] <= r_data[30530];
                
                r_data[30532] <= r_data[30531];
                
                r_data[30533] <= r_data[30532];
                
                r_data[30534] <= r_data[30533];
                
                r_data[30535] <= r_data[30534];
                
                r_data[30536] <= r_data[30535];
                
                r_data[30537] <= r_data[30536];
                
                r_data[30538] <= r_data[30537];
                
                r_data[30539] <= r_data[30538];
                
                r_data[30540] <= r_data[30539];
                
                r_data[30541] <= r_data[30540];
                
                r_data[30542] <= r_data[30541];
                
                r_data[30543] <= r_data[30542];
                
                r_data[30544] <= r_data[30543];
                
                r_data[30545] <= r_data[30544];
                
                r_data[30546] <= r_data[30545];
                
                r_data[30547] <= r_data[30546];
                
                r_data[30548] <= r_data[30547];
                
                r_data[30549] <= r_data[30548];
                
                r_data[30550] <= r_data[30549];
                
                r_data[30551] <= r_data[30550];
                
                r_data[30552] <= r_data[30551];
                
                r_data[30553] <= r_data[30552];
                
                r_data[30554] <= r_data[30553];
                
                r_data[30555] <= r_data[30554];
                
                r_data[30556] <= r_data[30555];
                
                r_data[30557] <= r_data[30556];
                
                r_data[30558] <= r_data[30557];
                
                r_data[30559] <= r_data[30558];
                
                r_data[30560] <= r_data[30559];
                
                r_data[30561] <= r_data[30560];
                
                r_data[30562] <= r_data[30561];
                
                r_data[30563] <= r_data[30562];
                
                r_data[30564] <= r_data[30563];
                
                r_data[30565] <= r_data[30564];
                
                r_data[30566] <= r_data[30565];
                
                r_data[30567] <= r_data[30566];
                
                r_data[30568] <= r_data[30567];
                
                r_data[30569] <= r_data[30568];
                
                r_data[30570] <= r_data[30569];
                
                r_data[30571] <= r_data[30570];
                
                r_data[30572] <= r_data[30571];
                
                r_data[30573] <= r_data[30572];
                
                r_data[30574] <= r_data[30573];
                
                r_data[30575] <= r_data[30574];
                
                r_data[30576] <= r_data[30575];
                
                r_data[30577] <= r_data[30576];
                
                r_data[30578] <= r_data[30577];
                
                r_data[30579] <= r_data[30578];
                
                r_data[30580] <= r_data[30579];
                
                r_data[30581] <= r_data[30580];
                
                r_data[30582] <= r_data[30581];
                
                r_data[30583] <= r_data[30582];
                
                r_data[30584] <= r_data[30583];
                
                r_data[30585] <= r_data[30584];
                
                r_data[30586] <= r_data[30585];
                
                r_data[30587] <= r_data[30586];
                
                r_data[30588] <= r_data[30587];
                
                r_data[30589] <= r_data[30588];
                
                r_data[30590] <= r_data[30589];
                
                r_data[30591] <= r_data[30590];
                
                r_data[30592] <= r_data[30591];
                
                r_data[30593] <= r_data[30592];
                
                r_data[30594] <= r_data[30593];
                
                r_data[30595] <= r_data[30594];
                
                r_data[30596] <= r_data[30595];
                
                r_data[30597] <= r_data[30596];
                
                r_data[30598] <= r_data[30597];
                
                r_data[30599] <= r_data[30598];
                
                r_data[30600] <= r_data[30599];
                
                r_data[30601] <= r_data[30600];
                
                r_data[30602] <= r_data[30601];
                
                r_data[30603] <= r_data[30602];
                
                r_data[30604] <= r_data[30603];
                
                r_data[30605] <= r_data[30604];
                
                r_data[30606] <= r_data[30605];
                
                r_data[30607] <= r_data[30606];
                
                r_data[30608] <= r_data[30607];
                
                r_data[30609] <= r_data[30608];
                
                r_data[30610] <= r_data[30609];
                
                r_data[30611] <= r_data[30610];
                
                r_data[30612] <= r_data[30611];
                
                r_data[30613] <= r_data[30612];
                
                r_data[30614] <= r_data[30613];
                
                r_data[30615] <= r_data[30614];
                
                r_data[30616] <= r_data[30615];
                
                r_data[30617] <= r_data[30616];
                
                r_data[30618] <= r_data[30617];
                
                r_data[30619] <= r_data[30618];
                
                r_data[30620] <= r_data[30619];
                
                r_data[30621] <= r_data[30620];
                
                r_data[30622] <= r_data[30621];
                
                r_data[30623] <= r_data[30622];
                
                r_data[30624] <= r_data[30623];
                
                r_data[30625] <= r_data[30624];
                
                r_data[30626] <= r_data[30625];
                
                r_data[30627] <= r_data[30626];
                
                r_data[30628] <= r_data[30627];
                
                r_data[30629] <= r_data[30628];
                
                r_data[30630] <= r_data[30629];
                
                r_data[30631] <= r_data[30630];
                
                r_data[30632] <= r_data[30631];
                
                r_data[30633] <= r_data[30632];
                
                r_data[30634] <= r_data[30633];
                
                r_data[30635] <= r_data[30634];
                
                r_data[30636] <= r_data[30635];
                
                r_data[30637] <= r_data[30636];
                
                r_data[30638] <= r_data[30637];
                
                r_data[30639] <= r_data[30638];
                
                r_data[30640] <= r_data[30639];
                
                r_data[30641] <= r_data[30640];
                
                r_data[30642] <= r_data[30641];
                
                r_data[30643] <= r_data[30642];
                
                r_data[30644] <= r_data[30643];
                
                r_data[30645] <= r_data[30644];
                
                r_data[30646] <= r_data[30645];
                
                r_data[30647] <= r_data[30646];
                
                r_data[30648] <= r_data[30647];
                
                r_data[30649] <= r_data[30648];
                
                r_data[30650] <= r_data[30649];
                
                r_data[30651] <= r_data[30650];
                
                r_data[30652] <= r_data[30651];
                
                r_data[30653] <= r_data[30652];
                
                r_data[30654] <= r_data[30653];
                
                r_data[30655] <= r_data[30654];
                
                r_data[30656] <= r_data[30655];
                
                r_data[30657] <= r_data[30656];
                
                r_data[30658] <= r_data[30657];
                
                r_data[30659] <= r_data[30658];
                
                r_data[30660] <= r_data[30659];
                
                r_data[30661] <= r_data[30660];
                
                r_data[30662] <= r_data[30661];
                
                r_data[30663] <= r_data[30662];
                
                r_data[30664] <= r_data[30663];
                
                r_data[30665] <= r_data[30664];
                
                r_data[30666] <= r_data[30665];
                
                r_data[30667] <= r_data[30666];
                
                r_data[30668] <= r_data[30667];
                
                r_data[30669] <= r_data[30668];
                
                r_data[30670] <= r_data[30669];
                
                r_data[30671] <= r_data[30670];
                
                r_data[30672] <= r_data[30671];
                
                r_data[30673] <= r_data[30672];
                
                r_data[30674] <= r_data[30673];
                
                r_data[30675] <= r_data[30674];
                
                r_data[30676] <= r_data[30675];
                
                r_data[30677] <= r_data[30676];
                
                r_data[30678] <= r_data[30677];
                
                r_data[30679] <= r_data[30678];
                
                r_data[30680] <= r_data[30679];
                
                r_data[30681] <= r_data[30680];
                
                r_data[30682] <= r_data[30681];
                
                r_data[30683] <= r_data[30682];
                
                r_data[30684] <= r_data[30683];
                
                r_data[30685] <= r_data[30684];
                
                r_data[30686] <= r_data[30685];
                
                r_data[30687] <= r_data[30686];
                
                r_data[30688] <= r_data[30687];
                
                r_data[30689] <= r_data[30688];
                
                r_data[30690] <= r_data[30689];
                
                r_data[30691] <= r_data[30690];
                
                r_data[30692] <= r_data[30691];
                
                r_data[30693] <= r_data[30692];
                
                r_data[30694] <= r_data[30693];
                
                r_data[30695] <= r_data[30694];
                
                r_data[30696] <= r_data[30695];
                
                r_data[30697] <= r_data[30696];
                
                r_data[30698] <= r_data[30697];
                
                r_data[30699] <= r_data[30698];
                
                r_data[30700] <= r_data[30699];
                
                r_data[30701] <= r_data[30700];
                
                r_data[30702] <= r_data[30701];
                
                r_data[30703] <= r_data[30702];
                
                r_data[30704] <= r_data[30703];
                
                r_data[30705] <= r_data[30704];
                
                r_data[30706] <= r_data[30705];
                
                r_data[30707] <= r_data[30706];
                
                r_data[30708] <= r_data[30707];
                
                r_data[30709] <= r_data[30708];
                
                r_data[30710] <= r_data[30709];
                
                r_data[30711] <= r_data[30710];
                
                r_data[30712] <= r_data[30711];
                
                r_data[30713] <= r_data[30712];
                
                r_data[30714] <= r_data[30713];
                
                r_data[30715] <= r_data[30714];
                
                r_data[30716] <= r_data[30715];
                
                r_data[30717] <= r_data[30716];
                
                r_data[30718] <= r_data[30717];
                
                r_data[30719] <= r_data[30718];
                
                r_data[30720] <= r_data[30719];
                
                r_data[30721] <= r_data[30720];
                
                r_data[30722] <= r_data[30721];
                
                r_data[30723] <= r_data[30722];
                
                r_data[30724] <= r_data[30723];
                
                r_data[30725] <= r_data[30724];
                
                r_data[30726] <= r_data[30725];
                
                r_data[30727] <= r_data[30726];
                
                r_data[30728] <= r_data[30727];
                
                r_data[30729] <= r_data[30728];
                
                r_data[30730] <= r_data[30729];
                
                r_data[30731] <= r_data[30730];
                
                r_data[30732] <= r_data[30731];
                
                r_data[30733] <= r_data[30732];
                
                r_data[30734] <= r_data[30733];
                
                r_data[30735] <= r_data[30734];
                
                r_data[30736] <= r_data[30735];
                
                r_data[30737] <= r_data[30736];
                
                r_data[30738] <= r_data[30737];
                
                r_data[30739] <= r_data[30738];
                
                r_data[30740] <= r_data[30739];
                
                r_data[30741] <= r_data[30740];
                
                r_data[30742] <= r_data[30741];
                
                r_data[30743] <= r_data[30742];
                
                r_data[30744] <= r_data[30743];
                
                r_data[30745] <= r_data[30744];
                
                r_data[30746] <= r_data[30745];
                
                r_data[30747] <= r_data[30746];
                
                r_data[30748] <= r_data[30747];
                
                r_data[30749] <= r_data[30748];
                
                r_data[30750] <= r_data[30749];
                
                r_data[30751] <= r_data[30750];
                
                r_data[30752] <= r_data[30751];
                
                r_data[30753] <= r_data[30752];
                
                r_data[30754] <= r_data[30753];
                
                r_data[30755] <= r_data[30754];
                
                r_data[30756] <= r_data[30755];
                
                r_data[30757] <= r_data[30756];
                
                r_data[30758] <= r_data[30757];
                
                r_data[30759] <= r_data[30758];
                
                r_data[30760] <= r_data[30759];
                
                r_data[30761] <= r_data[30760];
                
                r_data[30762] <= r_data[30761];
                
                r_data[30763] <= r_data[30762];
                
                r_data[30764] <= r_data[30763];
                
                r_data[30765] <= r_data[30764];
                
                r_data[30766] <= r_data[30765];
                
                r_data[30767] <= r_data[30766];
                
                r_data[30768] <= r_data[30767];
                
                r_data[30769] <= r_data[30768];
                
                r_data[30770] <= r_data[30769];
                
                r_data[30771] <= r_data[30770];
                
                r_data[30772] <= r_data[30771];
                
                r_data[30773] <= r_data[30772];
                
                r_data[30774] <= r_data[30773];
                
                r_data[30775] <= r_data[30774];
                
                r_data[30776] <= r_data[30775];
                
                r_data[30777] <= r_data[30776];
                
                r_data[30778] <= r_data[30777];
                
                r_data[30779] <= r_data[30778];
                
                r_data[30780] <= r_data[30779];
                
                r_data[30781] <= r_data[30780];
                
                r_data[30782] <= r_data[30781];
                
                r_data[30783] <= r_data[30782];
                
                r_data[30784] <= r_data[30783];
                
                r_data[30785] <= r_data[30784];
                
                r_data[30786] <= r_data[30785];
                
                r_data[30787] <= r_data[30786];
                
                r_data[30788] <= r_data[30787];
                
                r_data[30789] <= r_data[30788];
                
                r_data[30790] <= r_data[30789];
                
                r_data[30791] <= r_data[30790];
                
                r_data[30792] <= r_data[30791];
                
                r_data[30793] <= r_data[30792];
                
                r_data[30794] <= r_data[30793];
                
                r_data[30795] <= r_data[30794];
                
                r_data[30796] <= r_data[30795];
                
                r_data[30797] <= r_data[30796];
                
                r_data[30798] <= r_data[30797];
                
                r_data[30799] <= r_data[30798];
                
                r_data[30800] <= r_data[30799];
                
                r_data[30801] <= r_data[30800];
                
                r_data[30802] <= r_data[30801];
                
                r_data[30803] <= r_data[30802];
                
                r_data[30804] <= r_data[30803];
                
                r_data[30805] <= r_data[30804];
                
                r_data[30806] <= r_data[30805];
                
                r_data[30807] <= r_data[30806];
                
                r_data[30808] <= r_data[30807];
                
                r_data[30809] <= r_data[30808];
                
                r_data[30810] <= r_data[30809];
                
                r_data[30811] <= r_data[30810];
                
                r_data[30812] <= r_data[30811];
                
                r_data[30813] <= r_data[30812];
                
                r_data[30814] <= r_data[30813];
                
                r_data[30815] <= r_data[30814];
                
                r_data[30816] <= r_data[30815];
                
                r_data[30817] <= r_data[30816];
                
                r_data[30818] <= r_data[30817];
                
                r_data[30819] <= r_data[30818];
                
                r_data[30820] <= r_data[30819];
                
                r_data[30821] <= r_data[30820];
                
                r_data[30822] <= r_data[30821];
                
                r_data[30823] <= r_data[30822];
                
                r_data[30824] <= r_data[30823];
                
                r_data[30825] <= r_data[30824];
                
                r_data[30826] <= r_data[30825];
                
                r_data[30827] <= r_data[30826];
                
                r_data[30828] <= r_data[30827];
                
                r_data[30829] <= r_data[30828];
                
                r_data[30830] <= r_data[30829];
                
                r_data[30831] <= r_data[30830];
                
                r_data[30832] <= r_data[30831];
                
                r_data[30833] <= r_data[30832];
                
                r_data[30834] <= r_data[30833];
                
                r_data[30835] <= r_data[30834];
                
                r_data[30836] <= r_data[30835];
                
                r_data[30837] <= r_data[30836];
                
                r_data[30838] <= r_data[30837];
                
                r_data[30839] <= r_data[30838];
                
                r_data[30840] <= r_data[30839];
                
                r_data[30841] <= r_data[30840];
                
                r_data[30842] <= r_data[30841];
                
                r_data[30843] <= r_data[30842];
                
                r_data[30844] <= r_data[30843];
                
                r_data[30845] <= r_data[30844];
                
                r_data[30846] <= r_data[30845];
                
                r_data[30847] <= r_data[30846];
                
                r_data[30848] <= r_data[30847];
                
                r_data[30849] <= r_data[30848];
                
                r_data[30850] <= r_data[30849];
                
                r_data[30851] <= r_data[30850];
                
                r_data[30852] <= r_data[30851];
                
                r_data[30853] <= r_data[30852];
                
                r_data[30854] <= r_data[30853];
                
                r_data[30855] <= r_data[30854];
                
                r_data[30856] <= r_data[30855];
                
                r_data[30857] <= r_data[30856];
                
                r_data[30858] <= r_data[30857];
                
                r_data[30859] <= r_data[30858];
                
                r_data[30860] <= r_data[30859];
                
                r_data[30861] <= r_data[30860];
                
                r_data[30862] <= r_data[30861];
                
                r_data[30863] <= r_data[30862];
                
                r_data[30864] <= r_data[30863];
                
                r_data[30865] <= r_data[30864];
                
                r_data[30866] <= r_data[30865];
                
                r_data[30867] <= r_data[30866];
                
                r_data[30868] <= r_data[30867];
                
                r_data[30869] <= r_data[30868];
                
                r_data[30870] <= r_data[30869];
                
                r_data[30871] <= r_data[30870];
                
                r_data[30872] <= r_data[30871];
                
                r_data[30873] <= r_data[30872];
                
                r_data[30874] <= r_data[30873];
                
                r_data[30875] <= r_data[30874];
                
                r_data[30876] <= r_data[30875];
                
                r_data[30877] <= r_data[30876];
                
                r_data[30878] <= r_data[30877];
                
                r_data[30879] <= r_data[30878];
                
                r_data[30880] <= r_data[30879];
                
                r_data[30881] <= r_data[30880];
                
                r_data[30882] <= r_data[30881];
                
                r_data[30883] <= r_data[30882];
                
                r_data[30884] <= r_data[30883];
                
                r_data[30885] <= r_data[30884];
                
                r_data[30886] <= r_data[30885];
                
                r_data[30887] <= r_data[30886];
                
                r_data[30888] <= r_data[30887];
                
                r_data[30889] <= r_data[30888];
                
                r_data[30890] <= r_data[30889];
                
                r_data[30891] <= r_data[30890];
                
                r_data[30892] <= r_data[30891];
                
                r_data[30893] <= r_data[30892];
                
                r_data[30894] <= r_data[30893];
                
                r_data[30895] <= r_data[30894];
                
                r_data[30896] <= r_data[30895];
                
                r_data[30897] <= r_data[30896];
                
                r_data[30898] <= r_data[30897];
                
                r_data[30899] <= r_data[30898];
                
                r_data[30900] <= r_data[30899];
                
                r_data[30901] <= r_data[30900];
                
                r_data[30902] <= r_data[30901];
                
                r_data[30903] <= r_data[30902];
                
                r_data[30904] <= r_data[30903];
                
                r_data[30905] <= r_data[30904];
                
                r_data[30906] <= r_data[30905];
                
                r_data[30907] <= r_data[30906];
                
                r_data[30908] <= r_data[30907];
                
                r_data[30909] <= r_data[30908];
                
                r_data[30910] <= r_data[30909];
                
                r_data[30911] <= r_data[30910];
                
                r_data[30912] <= r_data[30911];
                
                r_data[30913] <= r_data[30912];
                
                r_data[30914] <= r_data[30913];
                
                r_data[30915] <= r_data[30914];
                
                r_data[30916] <= r_data[30915];
                
                r_data[30917] <= r_data[30916];
                
                r_data[30918] <= r_data[30917];
                
                r_data[30919] <= r_data[30918];
                
                r_data[30920] <= r_data[30919];
                
                r_data[30921] <= r_data[30920];
                
                r_data[30922] <= r_data[30921];
                
                r_data[30923] <= r_data[30922];
                
                r_data[30924] <= r_data[30923];
                
                r_data[30925] <= r_data[30924];
                
                r_data[30926] <= r_data[30925];
                
                r_data[30927] <= r_data[30926];
                
                r_data[30928] <= r_data[30927];
                
                r_data[30929] <= r_data[30928];
                
                r_data[30930] <= r_data[30929];
                
                r_data[30931] <= r_data[30930];
                
                r_data[30932] <= r_data[30931];
                
                r_data[30933] <= r_data[30932];
                
                r_data[30934] <= r_data[30933];
                
                r_data[30935] <= r_data[30934];
                
                r_data[30936] <= r_data[30935];
                
                r_data[30937] <= r_data[30936];
                
                r_data[30938] <= r_data[30937];
                
                r_data[30939] <= r_data[30938];
                
                r_data[30940] <= r_data[30939];
                
                r_data[30941] <= r_data[30940];
                
                r_data[30942] <= r_data[30941];
                
                r_data[30943] <= r_data[30942];
                
                r_data[30944] <= r_data[30943];
                
                r_data[30945] <= r_data[30944];
                
                r_data[30946] <= r_data[30945];
                
                r_data[30947] <= r_data[30946];
                
                r_data[30948] <= r_data[30947];
                
                r_data[30949] <= r_data[30948];
                
                r_data[30950] <= r_data[30949];
                
                r_data[30951] <= r_data[30950];
                
                r_data[30952] <= r_data[30951];
                
                r_data[30953] <= r_data[30952];
                
                r_data[30954] <= r_data[30953];
                
                r_data[30955] <= r_data[30954];
                
                r_data[30956] <= r_data[30955];
                
                r_data[30957] <= r_data[30956];
                
                r_data[30958] <= r_data[30957];
                
                r_data[30959] <= r_data[30958];
                
                r_data[30960] <= r_data[30959];
                
                r_data[30961] <= r_data[30960];
                
                r_data[30962] <= r_data[30961];
                
                r_data[30963] <= r_data[30962];
                
                r_data[30964] <= r_data[30963];
                
                r_data[30965] <= r_data[30964];
                
                r_data[30966] <= r_data[30965];
                
                r_data[30967] <= r_data[30966];
                
                r_data[30968] <= r_data[30967];
                
                r_data[30969] <= r_data[30968];
                
                r_data[30970] <= r_data[30969];
                
                r_data[30971] <= r_data[30970];
                
                r_data[30972] <= r_data[30971];
                
                r_data[30973] <= r_data[30972];
                
                r_data[30974] <= r_data[30973];
                
                r_data[30975] <= r_data[30974];
                
                r_data[30976] <= r_data[30975];
                
                r_data[30977] <= r_data[30976];
                
                r_data[30978] <= r_data[30977];
                
                r_data[30979] <= r_data[30978];
                
                r_data[30980] <= r_data[30979];
                
                r_data[30981] <= r_data[30980];
                
                r_data[30982] <= r_data[30981];
                
                r_data[30983] <= r_data[30982];
                
                r_data[30984] <= r_data[30983];
                
                r_data[30985] <= r_data[30984];
                
                r_data[30986] <= r_data[30985];
                
                r_data[30987] <= r_data[30986];
                
                r_data[30988] <= r_data[30987];
                
                r_data[30989] <= r_data[30988];
                
                r_data[30990] <= r_data[30989];
                
                r_data[30991] <= r_data[30990];
                
                r_data[30992] <= r_data[30991];
                
                r_data[30993] <= r_data[30992];
                
                r_data[30994] <= r_data[30993];
                
                r_data[30995] <= r_data[30994];
                
                r_data[30996] <= r_data[30995];
                
                r_data[30997] <= r_data[30996];
                
                r_data[30998] <= r_data[30997];
                
                r_data[30999] <= r_data[30998];
                
                r_data[31000] <= r_data[30999];
                
                r_data[31001] <= r_data[31000];
                
                r_data[31002] <= r_data[31001];
                
                r_data[31003] <= r_data[31002];
                
                r_data[31004] <= r_data[31003];
                
                r_data[31005] <= r_data[31004];
                
                r_data[31006] <= r_data[31005];
                
                r_data[31007] <= r_data[31006];
                
                r_data[31008] <= r_data[31007];
                
                r_data[31009] <= r_data[31008];
                
                r_data[31010] <= r_data[31009];
                
                r_data[31011] <= r_data[31010];
                
                r_data[31012] <= r_data[31011];
                
                r_data[31013] <= r_data[31012];
                
                r_data[31014] <= r_data[31013];
                
                r_data[31015] <= r_data[31014];
                
                r_data[31016] <= r_data[31015];
                
                r_data[31017] <= r_data[31016];
                
                r_data[31018] <= r_data[31017];
                
                r_data[31019] <= r_data[31018];
                
                r_data[31020] <= r_data[31019];
                
                r_data[31021] <= r_data[31020];
                
                r_data[31022] <= r_data[31021];
                
                r_data[31023] <= r_data[31022];
                
                r_data[31024] <= r_data[31023];
                
                r_data[31025] <= r_data[31024];
                
                r_data[31026] <= r_data[31025];
                
                r_data[31027] <= r_data[31026];
                
                r_data[31028] <= r_data[31027];
                
                r_data[31029] <= r_data[31028];
                
                r_data[31030] <= r_data[31029];
                
                r_data[31031] <= r_data[31030];
                
                r_data[31032] <= r_data[31031];
                
                r_data[31033] <= r_data[31032];
                
                r_data[31034] <= r_data[31033];
                
                r_data[31035] <= r_data[31034];
                
                r_data[31036] <= r_data[31035];
                
                r_data[31037] <= r_data[31036];
                
                r_data[31038] <= r_data[31037];
                
                r_data[31039] <= r_data[31038];
                
                r_data[31040] <= r_data[31039];
                
                r_data[31041] <= r_data[31040];
                
                r_data[31042] <= r_data[31041];
                
                r_data[31043] <= r_data[31042];
                
                r_data[31044] <= r_data[31043];
                
                r_data[31045] <= r_data[31044];
                
                r_data[31046] <= r_data[31045];
                
                r_data[31047] <= r_data[31046];
                
                r_data[31048] <= r_data[31047];
                
                r_data[31049] <= r_data[31048];
                
                r_data[31050] <= r_data[31049];
                
                r_data[31051] <= r_data[31050];
                
                r_data[31052] <= r_data[31051];
                
                r_data[31053] <= r_data[31052];
                
                r_data[31054] <= r_data[31053];
                
                r_data[31055] <= r_data[31054];
                
                r_data[31056] <= r_data[31055];
                
                r_data[31057] <= r_data[31056];
                
                r_data[31058] <= r_data[31057];
                
                r_data[31059] <= r_data[31058];
                
                r_data[31060] <= r_data[31059];
                
                r_data[31061] <= r_data[31060];
                
                r_data[31062] <= r_data[31061];
                
                r_data[31063] <= r_data[31062];
                
                r_data[31064] <= r_data[31063];
                
                r_data[31065] <= r_data[31064];
                
                r_data[31066] <= r_data[31065];
                
                r_data[31067] <= r_data[31066];
                
                r_data[31068] <= r_data[31067];
                
                r_data[31069] <= r_data[31068];
                
                r_data[31070] <= r_data[31069];
                
                r_data[31071] <= r_data[31070];
                
                r_data[31072] <= r_data[31071];
                
                r_data[31073] <= r_data[31072];
                
                r_data[31074] <= r_data[31073];
                
                r_data[31075] <= r_data[31074];
                
                r_data[31076] <= r_data[31075];
                
                r_data[31077] <= r_data[31076];
                
                r_data[31078] <= r_data[31077];
                
                r_data[31079] <= r_data[31078];
                
                r_data[31080] <= r_data[31079];
                
                r_data[31081] <= r_data[31080];
                
                r_data[31082] <= r_data[31081];
                
                r_data[31083] <= r_data[31082];
                
                r_data[31084] <= r_data[31083];
                
                r_data[31085] <= r_data[31084];
                
                r_data[31086] <= r_data[31085];
                
                r_data[31087] <= r_data[31086];
                
                r_data[31088] <= r_data[31087];
                
                r_data[31089] <= r_data[31088];
                
                r_data[31090] <= r_data[31089];
                
                r_data[31091] <= r_data[31090];
                
                r_data[31092] <= r_data[31091];
                
                r_data[31093] <= r_data[31092];
                
                r_data[31094] <= r_data[31093];
                
                r_data[31095] <= r_data[31094];
                
                r_data[31096] <= r_data[31095];
                
                r_data[31097] <= r_data[31096];
                
                r_data[31098] <= r_data[31097];
                
                r_data[31099] <= r_data[31098];
                
                r_data[31100] <= r_data[31099];
                
                r_data[31101] <= r_data[31100];
                
                r_data[31102] <= r_data[31101];
                
                r_data[31103] <= r_data[31102];
                
                r_data[31104] <= r_data[31103];
                
                r_data[31105] <= r_data[31104];
                
                r_data[31106] <= r_data[31105];
                
                r_data[31107] <= r_data[31106];
                
                r_data[31108] <= r_data[31107];
                
                r_data[31109] <= r_data[31108];
                
                r_data[31110] <= r_data[31109];
                
                r_data[31111] <= r_data[31110];
                
                r_data[31112] <= r_data[31111];
                
                r_data[31113] <= r_data[31112];
                
                r_data[31114] <= r_data[31113];
                
                r_data[31115] <= r_data[31114];
                
                r_data[31116] <= r_data[31115];
                
                r_data[31117] <= r_data[31116];
                
                r_data[31118] <= r_data[31117];
                
                r_data[31119] <= r_data[31118];
                
                r_data[31120] <= r_data[31119];
                
                r_data[31121] <= r_data[31120];
                
                r_data[31122] <= r_data[31121];
                
                r_data[31123] <= r_data[31122];
                
                r_data[31124] <= r_data[31123];
                
                r_data[31125] <= r_data[31124];
                
                r_data[31126] <= r_data[31125];
                
                r_data[31127] <= r_data[31126];
                
                r_data[31128] <= r_data[31127];
                
                r_data[31129] <= r_data[31128];
                
                r_data[31130] <= r_data[31129];
                
                r_data[31131] <= r_data[31130];
                
                r_data[31132] <= r_data[31131];
                
                r_data[31133] <= r_data[31132];
                
                r_data[31134] <= r_data[31133];
                
                r_data[31135] <= r_data[31134];
                
                r_data[31136] <= r_data[31135];
                
                r_data[31137] <= r_data[31136];
                
                r_data[31138] <= r_data[31137];
                
                r_data[31139] <= r_data[31138];
                
                r_data[31140] <= r_data[31139];
                
                r_data[31141] <= r_data[31140];
                
                r_data[31142] <= r_data[31141];
                
                r_data[31143] <= r_data[31142];
                
                r_data[31144] <= r_data[31143];
                
                r_data[31145] <= r_data[31144];
                
                r_data[31146] <= r_data[31145];
                
                r_data[31147] <= r_data[31146];
                
                r_data[31148] <= r_data[31147];
                
                r_data[31149] <= r_data[31148];
                
                r_data[31150] <= r_data[31149];
                
                r_data[31151] <= r_data[31150];
                
                r_data[31152] <= r_data[31151];
                
                r_data[31153] <= r_data[31152];
                
                r_data[31154] <= r_data[31153];
                
                r_data[31155] <= r_data[31154];
                
                r_data[31156] <= r_data[31155];
                
                r_data[31157] <= r_data[31156];
                
                r_data[31158] <= r_data[31157];
                
                r_data[31159] <= r_data[31158];
                
                r_data[31160] <= r_data[31159];
                
                r_data[31161] <= r_data[31160];
                
                r_data[31162] <= r_data[31161];
                
                r_data[31163] <= r_data[31162];
                
                r_data[31164] <= r_data[31163];
                
                r_data[31165] <= r_data[31164];
                
                r_data[31166] <= r_data[31165];
                
                r_data[31167] <= r_data[31166];
                
                r_data[31168] <= r_data[31167];
                
                r_data[31169] <= r_data[31168];
                
                r_data[31170] <= r_data[31169];
                
                r_data[31171] <= r_data[31170];
                
                r_data[31172] <= r_data[31171];
                
                r_data[31173] <= r_data[31172];
                
                r_data[31174] <= r_data[31173];
                
                r_data[31175] <= r_data[31174];
                
                r_data[31176] <= r_data[31175];
                
                r_data[31177] <= r_data[31176];
                
                r_data[31178] <= r_data[31177];
                
                r_data[31179] <= r_data[31178];
                
                r_data[31180] <= r_data[31179];
                
                r_data[31181] <= r_data[31180];
                
                r_data[31182] <= r_data[31181];
                
                r_data[31183] <= r_data[31182];
                
                r_data[31184] <= r_data[31183];
                
                r_data[31185] <= r_data[31184];
                
                r_data[31186] <= r_data[31185];
                
                r_data[31187] <= r_data[31186];
                
                r_data[31188] <= r_data[31187];
                
                r_data[31189] <= r_data[31188];
                
                r_data[31190] <= r_data[31189];
                
                r_data[31191] <= r_data[31190];
                
                r_data[31192] <= r_data[31191];
                
                r_data[31193] <= r_data[31192];
                
                r_data[31194] <= r_data[31193];
                
                r_data[31195] <= r_data[31194];
                
                r_data[31196] <= r_data[31195];
                
                r_data[31197] <= r_data[31196];
                
                r_data[31198] <= r_data[31197];
                
                r_data[31199] <= r_data[31198];
                
                r_data[31200] <= r_data[31199];
                
                r_data[31201] <= r_data[31200];
                
                r_data[31202] <= r_data[31201];
                
                r_data[31203] <= r_data[31202];
                
                r_data[31204] <= r_data[31203];
                
                r_data[31205] <= r_data[31204];
                
                r_data[31206] <= r_data[31205];
                
                r_data[31207] <= r_data[31206];
                
                r_data[31208] <= r_data[31207];
                
                r_data[31209] <= r_data[31208];
                
                r_data[31210] <= r_data[31209];
                
                r_data[31211] <= r_data[31210];
                
                r_data[31212] <= r_data[31211];
                
                r_data[31213] <= r_data[31212];
                
                r_data[31214] <= r_data[31213];
                
                r_data[31215] <= r_data[31214];
                
                r_data[31216] <= r_data[31215];
                
                r_data[31217] <= r_data[31216];
                
                r_data[31218] <= r_data[31217];
                
                r_data[31219] <= r_data[31218];
                
                r_data[31220] <= r_data[31219];
                
                r_data[31221] <= r_data[31220];
                
                r_data[31222] <= r_data[31221];
                
                r_data[31223] <= r_data[31222];
                
                r_data[31224] <= r_data[31223];
                
                r_data[31225] <= r_data[31224];
                
                r_data[31226] <= r_data[31225];
                
                r_data[31227] <= r_data[31226];
                
                r_data[31228] <= r_data[31227];
                
                r_data[31229] <= r_data[31228];
                
                r_data[31230] <= r_data[31229];
                
                r_data[31231] <= r_data[31230];
                
                r_data[31232] <= r_data[31231];
                
                r_data[31233] <= r_data[31232];
                
                r_data[31234] <= r_data[31233];
                
                r_data[31235] <= r_data[31234];
                
                r_data[31236] <= r_data[31235];
                
                r_data[31237] <= r_data[31236];
                
                r_data[31238] <= r_data[31237];
                
                r_data[31239] <= r_data[31238];
                
                r_data[31240] <= r_data[31239];
                
                r_data[31241] <= r_data[31240];
                
                r_data[31242] <= r_data[31241];
                
                r_data[31243] <= r_data[31242];
                
                r_data[31244] <= r_data[31243];
                
                r_data[31245] <= r_data[31244];
                
                r_data[31246] <= r_data[31245];
                
                r_data[31247] <= r_data[31246];
                
                r_data[31248] <= r_data[31247];
                
                r_data[31249] <= r_data[31248];
                
                r_data[31250] <= r_data[31249];
                
                r_data[31251] <= r_data[31250];
                
                r_data[31252] <= r_data[31251];
                
                r_data[31253] <= r_data[31252];
                
                r_data[31254] <= r_data[31253];
                
                r_data[31255] <= r_data[31254];
                
                r_data[31256] <= r_data[31255];
                
                r_data[31257] <= r_data[31256];
                
                r_data[31258] <= r_data[31257];
                
                r_data[31259] <= r_data[31258];
                
                r_data[31260] <= r_data[31259];
                
                r_data[31261] <= r_data[31260];
                
                r_data[31262] <= r_data[31261];
                
                r_data[31263] <= r_data[31262];
                
                r_data[31264] <= r_data[31263];
                
                r_data[31265] <= r_data[31264];
                
                r_data[31266] <= r_data[31265];
                
                r_data[31267] <= r_data[31266];
                
                r_data[31268] <= r_data[31267];
                
                r_data[31269] <= r_data[31268];
                
                r_data[31270] <= r_data[31269];
                
                r_data[31271] <= r_data[31270];
                
                r_data[31272] <= r_data[31271];
                
                r_data[31273] <= r_data[31272];
                
                r_data[31274] <= r_data[31273];
                
                r_data[31275] <= r_data[31274];
                
                r_data[31276] <= r_data[31275];
                
                r_data[31277] <= r_data[31276];
                
                r_data[31278] <= r_data[31277];
                
                r_data[31279] <= r_data[31278];
                
                r_data[31280] <= r_data[31279];
                
                r_data[31281] <= r_data[31280];
                
                r_data[31282] <= r_data[31281];
                
                r_data[31283] <= r_data[31282];
                
                r_data[31284] <= r_data[31283];
                
                r_data[31285] <= r_data[31284];
                
                r_data[31286] <= r_data[31285];
                
                r_data[31287] <= r_data[31286];
                
                r_data[31288] <= r_data[31287];
                
                r_data[31289] <= r_data[31288];
                
                r_data[31290] <= r_data[31289];
                
                r_data[31291] <= r_data[31290];
                
                r_data[31292] <= r_data[31291];
                
                r_data[31293] <= r_data[31292];
                
                r_data[31294] <= r_data[31293];
                
                r_data[31295] <= r_data[31294];
                
                r_data[31296] <= r_data[31295];
                
                r_data[31297] <= r_data[31296];
                
                r_data[31298] <= r_data[31297];
                
                r_data[31299] <= r_data[31298];
                
                r_data[31300] <= r_data[31299];
                
                r_data[31301] <= r_data[31300];
                
                r_data[31302] <= r_data[31301];
                
                r_data[31303] <= r_data[31302];
                
                r_data[31304] <= r_data[31303];
                
                r_data[31305] <= r_data[31304];
                
                r_data[31306] <= r_data[31305];
                
                r_data[31307] <= r_data[31306];
                
                r_data[31308] <= r_data[31307];
                
                r_data[31309] <= r_data[31308];
                
                r_data[31310] <= r_data[31309];
                
                r_data[31311] <= r_data[31310];
                
                r_data[31312] <= r_data[31311];
                
                r_data[31313] <= r_data[31312];
                
                r_data[31314] <= r_data[31313];
                
                r_data[31315] <= r_data[31314];
                
                r_data[31316] <= r_data[31315];
                
                r_data[31317] <= r_data[31316];
                
                r_data[31318] <= r_data[31317];
                
                r_data[31319] <= r_data[31318];
                
                r_data[31320] <= r_data[31319];
                
                r_data[31321] <= r_data[31320];
                
                r_data[31322] <= r_data[31321];
                
                r_data[31323] <= r_data[31322];
                
                r_data[31324] <= r_data[31323];
                
                r_data[31325] <= r_data[31324];
                
                r_data[31326] <= r_data[31325];
                
                r_data[31327] <= r_data[31326];
                
                r_data[31328] <= r_data[31327];
                
                r_data[31329] <= r_data[31328];
                
                r_data[31330] <= r_data[31329];
                
                r_data[31331] <= r_data[31330];
                
                r_data[31332] <= r_data[31331];
                
                r_data[31333] <= r_data[31332];
                
                r_data[31334] <= r_data[31333];
                
                r_data[31335] <= r_data[31334];
                
                r_data[31336] <= r_data[31335];
                
                r_data[31337] <= r_data[31336];
                
                r_data[31338] <= r_data[31337];
                
                r_data[31339] <= r_data[31338];
                
                r_data[31340] <= r_data[31339];
                
                r_data[31341] <= r_data[31340];
                
                r_data[31342] <= r_data[31341];
                
                r_data[31343] <= r_data[31342];
                
                r_data[31344] <= r_data[31343];
                
                r_data[31345] <= r_data[31344];
                
                r_data[31346] <= r_data[31345];
                
                r_data[31347] <= r_data[31346];
                
                r_data[31348] <= r_data[31347];
                
                r_data[31349] <= r_data[31348];
                
                r_data[31350] <= r_data[31349];
                
                r_data[31351] <= r_data[31350];
                
                r_data[31352] <= r_data[31351];
                
                r_data[31353] <= r_data[31352];
                
                r_data[31354] <= r_data[31353];
                
                r_data[31355] <= r_data[31354];
                
                r_data[31356] <= r_data[31355];
                
                r_data[31357] <= r_data[31356];
                
                r_data[31358] <= r_data[31357];
                
                r_data[31359] <= r_data[31358];
                
                r_data[31360] <= r_data[31359];
                
                r_data[31361] <= r_data[31360];
                
                r_data[31362] <= r_data[31361];
                
                r_data[31363] <= r_data[31362];
                
                r_data[31364] <= r_data[31363];
                
                r_data[31365] <= r_data[31364];
                
                r_data[31366] <= r_data[31365];
                
                r_data[31367] <= r_data[31366];
                
                r_data[31368] <= r_data[31367];
                
                r_data[31369] <= r_data[31368];
                
                r_data[31370] <= r_data[31369];
                
                r_data[31371] <= r_data[31370];
                
                r_data[31372] <= r_data[31371];
                
                r_data[31373] <= r_data[31372];
                
                r_data[31374] <= r_data[31373];
                
                r_data[31375] <= r_data[31374];
                
                r_data[31376] <= r_data[31375];
                
                r_data[31377] <= r_data[31376];
                
                r_data[31378] <= r_data[31377];
                
                r_data[31379] <= r_data[31378];
                
                r_data[31380] <= r_data[31379];
                
                r_data[31381] <= r_data[31380];
                
                r_data[31382] <= r_data[31381];
                
                r_data[31383] <= r_data[31382];
                
                r_data[31384] <= r_data[31383];
                
                r_data[31385] <= r_data[31384];
                
                r_data[31386] <= r_data[31385];
                
                r_data[31387] <= r_data[31386];
                
                r_data[31388] <= r_data[31387];
                
                r_data[31389] <= r_data[31388];
                
                r_data[31390] <= r_data[31389];
                
                r_data[31391] <= r_data[31390];
                
                r_data[31392] <= r_data[31391];
                
                r_data[31393] <= r_data[31392];
                
                r_data[31394] <= r_data[31393];
                
                r_data[31395] <= r_data[31394];
                
                r_data[31396] <= r_data[31395];
                
                r_data[31397] <= r_data[31396];
                
                r_data[31398] <= r_data[31397];
                
                r_data[31399] <= r_data[31398];
                
                r_data[31400] <= r_data[31399];
                
                r_data[31401] <= r_data[31400];
                
                r_data[31402] <= r_data[31401];
                
                r_data[31403] <= r_data[31402];
                
                r_data[31404] <= r_data[31403];
                
                r_data[31405] <= r_data[31404];
                
                r_data[31406] <= r_data[31405];
                
                r_data[31407] <= r_data[31406];
                
                r_data[31408] <= r_data[31407];
                
                r_data[31409] <= r_data[31408];
                
                r_data[31410] <= r_data[31409];
                
                r_data[31411] <= r_data[31410];
                
                r_data[31412] <= r_data[31411];
                
                r_data[31413] <= r_data[31412];
                
                r_data[31414] <= r_data[31413];
                
                r_data[31415] <= r_data[31414];
                
                r_data[31416] <= r_data[31415];
                
                r_data[31417] <= r_data[31416];
                
                r_data[31418] <= r_data[31417];
                
                r_data[31419] <= r_data[31418];
                
                r_data[31420] <= r_data[31419];
                
                r_data[31421] <= r_data[31420];
                
                r_data[31422] <= r_data[31421];
                
                r_data[31423] <= r_data[31422];
                
                r_data[31424] <= r_data[31423];
                
                r_data[31425] <= r_data[31424];
                
                r_data[31426] <= r_data[31425];
                
                r_data[31427] <= r_data[31426];
                
                r_data[31428] <= r_data[31427];
                
                r_data[31429] <= r_data[31428];
                
                r_data[31430] <= r_data[31429];
                
                r_data[31431] <= r_data[31430];
                
                r_data[31432] <= r_data[31431];
                
                r_data[31433] <= r_data[31432];
                
                r_data[31434] <= r_data[31433];
                
                r_data[31435] <= r_data[31434];
                
                r_data[31436] <= r_data[31435];
                
                r_data[31437] <= r_data[31436];
                
                r_data[31438] <= r_data[31437];
                
                r_data[31439] <= r_data[31438];
                
                r_data[31440] <= r_data[31439];
                
                r_data[31441] <= r_data[31440];
                
                r_data[31442] <= r_data[31441];
                
                r_data[31443] <= r_data[31442];
                
                r_data[31444] <= r_data[31443];
                
                r_data[31445] <= r_data[31444];
                
                r_data[31446] <= r_data[31445];
                
                r_data[31447] <= r_data[31446];
                
                r_data[31448] <= r_data[31447];
                
                r_data[31449] <= r_data[31448];
                
                r_data[31450] <= r_data[31449];
                
                r_data[31451] <= r_data[31450];
                
                r_data[31452] <= r_data[31451];
                
                r_data[31453] <= r_data[31452];
                
                r_data[31454] <= r_data[31453];
                
                r_data[31455] <= r_data[31454];
                
                r_data[31456] <= r_data[31455];
                
                r_data[31457] <= r_data[31456];
                
                r_data[31458] <= r_data[31457];
                
                r_data[31459] <= r_data[31458];
                
                r_data[31460] <= r_data[31459];
                
                r_data[31461] <= r_data[31460];
                
                r_data[31462] <= r_data[31461];
                
                r_data[31463] <= r_data[31462];
                
                r_data[31464] <= r_data[31463];
                
                r_data[31465] <= r_data[31464];
                
                r_data[31466] <= r_data[31465];
                
                r_data[31467] <= r_data[31466];
                
                r_data[31468] <= r_data[31467];
                
                r_data[31469] <= r_data[31468];
                
                r_data[31470] <= r_data[31469];
                
                r_data[31471] <= r_data[31470];
                
                r_data[31472] <= r_data[31471];
                
                r_data[31473] <= r_data[31472];
                
                r_data[31474] <= r_data[31473];
                
                r_data[31475] <= r_data[31474];
                
                r_data[31476] <= r_data[31475];
                
                r_data[31477] <= r_data[31476];
                
                r_data[31478] <= r_data[31477];
                
                r_data[31479] <= r_data[31478];
                
                r_data[31480] <= r_data[31479];
                
                r_data[31481] <= r_data[31480];
                
                r_data[31482] <= r_data[31481];
                
                r_data[31483] <= r_data[31482];
                
                r_data[31484] <= r_data[31483];
                
                r_data[31485] <= r_data[31484];
                
                r_data[31486] <= r_data[31485];
                
                r_data[31487] <= r_data[31486];
                
                r_data[31488] <= r_data[31487];
                
                r_data[31489] <= r_data[31488];
                
                r_data[31490] <= r_data[31489];
                
                r_data[31491] <= r_data[31490];
                
                r_data[31492] <= r_data[31491];
                
                r_data[31493] <= r_data[31492];
                
                r_data[31494] <= r_data[31493];
                
                r_data[31495] <= r_data[31494];
                
                r_data[31496] <= r_data[31495];
                
                r_data[31497] <= r_data[31496];
                
                r_data[31498] <= r_data[31497];
                
                r_data[31499] <= r_data[31498];
                
                r_data[31500] <= r_data[31499];
                
                r_data[31501] <= r_data[31500];
                
                r_data[31502] <= r_data[31501];
                
                r_data[31503] <= r_data[31502];
                
                r_data[31504] <= r_data[31503];
                
                r_data[31505] <= r_data[31504];
                
                r_data[31506] <= r_data[31505];
                
                r_data[31507] <= r_data[31506];
                
                r_data[31508] <= r_data[31507];
                
                r_data[31509] <= r_data[31508];
                
                r_data[31510] <= r_data[31509];
                
                r_data[31511] <= r_data[31510];
                
                r_data[31512] <= r_data[31511];
                
                r_data[31513] <= r_data[31512];
                
                r_data[31514] <= r_data[31513];
                
                r_data[31515] <= r_data[31514];
                
                r_data[31516] <= r_data[31515];
                
                r_data[31517] <= r_data[31516];
                
                r_data[31518] <= r_data[31517];
                
                r_data[31519] <= r_data[31518];
                
                r_data[31520] <= r_data[31519];
                
                r_data[31521] <= r_data[31520];
                
                r_data[31522] <= r_data[31521];
                
                r_data[31523] <= r_data[31522];
                
                r_data[31524] <= r_data[31523];
                
                r_data[31525] <= r_data[31524];
                
                r_data[31526] <= r_data[31525];
                
                r_data[31527] <= r_data[31526];
                
                r_data[31528] <= r_data[31527];
                
                r_data[31529] <= r_data[31528];
                
                r_data[31530] <= r_data[31529];
                
                r_data[31531] <= r_data[31530];
                
                r_data[31532] <= r_data[31531];
                
                r_data[31533] <= r_data[31532];
                
                r_data[31534] <= r_data[31533];
                
                r_data[31535] <= r_data[31534];
                
                r_data[31536] <= r_data[31535];
                
                r_data[31537] <= r_data[31536];
                
                r_data[31538] <= r_data[31537];
                
                r_data[31539] <= r_data[31538];
                
                r_data[31540] <= r_data[31539];
                
                r_data[31541] <= r_data[31540];
                
                r_data[31542] <= r_data[31541];
                
                r_data[31543] <= r_data[31542];
                
                r_data[31544] <= r_data[31543];
                
                r_data[31545] <= r_data[31544];
                
                r_data[31546] <= r_data[31545];
                
                r_data[31547] <= r_data[31546];
                
                r_data[31548] <= r_data[31547];
                
                r_data[31549] <= r_data[31548];
                
                r_data[31550] <= r_data[31549];
                
                r_data[31551] <= r_data[31550];
                
                r_data[31552] <= r_data[31551];
                
                r_data[31553] <= r_data[31552];
                
                r_data[31554] <= r_data[31553];
                
                r_data[31555] <= r_data[31554];
                
                r_data[31556] <= r_data[31555];
                
                r_data[31557] <= r_data[31556];
                
                r_data[31558] <= r_data[31557];
                
                r_data[31559] <= r_data[31558];
                
                r_data[31560] <= r_data[31559];
                
                r_data[31561] <= r_data[31560];
                
                r_data[31562] <= r_data[31561];
                
                r_data[31563] <= r_data[31562];
                
                r_data[31564] <= r_data[31563];
                
                r_data[31565] <= r_data[31564];
                
                r_data[31566] <= r_data[31565];
                
                r_data[31567] <= r_data[31566];
                
                r_data[31568] <= r_data[31567];
                
                r_data[31569] <= r_data[31568];
                
                r_data[31570] <= r_data[31569];
                
                r_data[31571] <= r_data[31570];
                
                r_data[31572] <= r_data[31571];
                
                r_data[31573] <= r_data[31572];
                
                r_data[31574] <= r_data[31573];
                
                r_data[31575] <= r_data[31574];
                
                r_data[31576] <= r_data[31575];
                
                r_data[31577] <= r_data[31576];
                
                r_data[31578] <= r_data[31577];
                
                r_data[31579] <= r_data[31578];
                
                r_data[31580] <= r_data[31579];
                
                r_data[31581] <= r_data[31580];
                
                r_data[31582] <= r_data[31581];
                
                r_data[31583] <= r_data[31582];
                
                r_data[31584] <= r_data[31583];
                
                r_data[31585] <= r_data[31584];
                
                r_data[31586] <= r_data[31585];
                
                r_data[31587] <= r_data[31586];
                
                r_data[31588] <= r_data[31587];
                
                r_data[31589] <= r_data[31588];
                
                r_data[31590] <= r_data[31589];
                
                r_data[31591] <= r_data[31590];
                
                r_data[31592] <= r_data[31591];
                
                r_data[31593] <= r_data[31592];
                
                r_data[31594] <= r_data[31593];
                
                r_data[31595] <= r_data[31594];
                
                r_data[31596] <= r_data[31595];
                
                r_data[31597] <= r_data[31596];
                
                r_data[31598] <= r_data[31597];
                
                r_data[31599] <= r_data[31598];
                
                r_data[31600] <= r_data[31599];
                
                r_data[31601] <= r_data[31600];
                
                r_data[31602] <= r_data[31601];
                
                r_data[31603] <= r_data[31602];
                
                r_data[31604] <= r_data[31603];
                
                r_data[31605] <= r_data[31604];
                
                r_data[31606] <= r_data[31605];
                
                r_data[31607] <= r_data[31606];
                
                r_data[31608] <= r_data[31607];
                
                r_data[31609] <= r_data[31608];
                
                r_data[31610] <= r_data[31609];
                
                r_data[31611] <= r_data[31610];
                
                r_data[31612] <= r_data[31611];
                
                r_data[31613] <= r_data[31612];
                
                r_data[31614] <= r_data[31613];
                
                r_data[31615] <= r_data[31614];
                
                r_data[31616] <= r_data[31615];
                
                r_data[31617] <= r_data[31616];
                
                r_data[31618] <= r_data[31617];
                
                r_data[31619] <= r_data[31618];
                
                r_data[31620] <= r_data[31619];
                
                r_data[31621] <= r_data[31620];
                
                r_data[31622] <= r_data[31621];
                
                r_data[31623] <= r_data[31622];
                
                r_data[31624] <= r_data[31623];
                
                r_data[31625] <= r_data[31624];
                
                r_data[31626] <= r_data[31625];
                
                r_data[31627] <= r_data[31626];
                
                r_data[31628] <= r_data[31627];
                
                r_data[31629] <= r_data[31628];
                
                r_data[31630] <= r_data[31629];
                
                r_data[31631] <= r_data[31630];
                
                r_data[31632] <= r_data[31631];
                
                r_data[31633] <= r_data[31632];
                
                r_data[31634] <= r_data[31633];
                
                r_data[31635] <= r_data[31634];
                
                r_data[31636] <= r_data[31635];
                
                r_data[31637] <= r_data[31636];
                
                r_data[31638] <= r_data[31637];
                
                r_data[31639] <= r_data[31638];
                
                r_data[31640] <= r_data[31639];
                
                r_data[31641] <= r_data[31640];
                
                r_data[31642] <= r_data[31641];
                
                r_data[31643] <= r_data[31642];
                
                r_data[31644] <= r_data[31643];
                
                r_data[31645] <= r_data[31644];
                
                r_data[31646] <= r_data[31645];
                
                r_data[31647] <= r_data[31646];
                
                r_data[31648] <= r_data[31647];
                
                r_data[31649] <= r_data[31648];
                
                r_data[31650] <= r_data[31649];
                
                r_data[31651] <= r_data[31650];
                
                r_data[31652] <= r_data[31651];
                
                r_data[31653] <= r_data[31652];
                
                r_data[31654] <= r_data[31653];
                
                r_data[31655] <= r_data[31654];
                
                r_data[31656] <= r_data[31655];
                
                r_data[31657] <= r_data[31656];
                
                r_data[31658] <= r_data[31657];
                
                r_data[31659] <= r_data[31658];
                
                r_data[31660] <= r_data[31659];
                
                r_data[31661] <= r_data[31660];
                
                r_data[31662] <= r_data[31661];
                
                r_data[31663] <= r_data[31662];
                
                r_data[31664] <= r_data[31663];
                
                r_data[31665] <= r_data[31664];
                
                r_data[31666] <= r_data[31665];
                
                r_data[31667] <= r_data[31666];
                
                r_data[31668] <= r_data[31667];
                
                r_data[31669] <= r_data[31668];
                
                r_data[31670] <= r_data[31669];
                
                r_data[31671] <= r_data[31670];
                
                r_data[31672] <= r_data[31671];
                
                r_data[31673] <= r_data[31672];
                
                r_data[31674] <= r_data[31673];
                
                r_data[31675] <= r_data[31674];
                
                r_data[31676] <= r_data[31675];
                
                r_data[31677] <= r_data[31676];
                
                r_data[31678] <= r_data[31677];
                
                r_data[31679] <= r_data[31678];
                
                r_data[31680] <= r_data[31679];
                
                r_data[31681] <= r_data[31680];
                
                r_data[31682] <= r_data[31681];
                
                r_data[31683] <= r_data[31682];
                
                r_data[31684] <= r_data[31683];
                
                r_data[31685] <= r_data[31684];
                
                r_data[31686] <= r_data[31685];
                
                r_data[31687] <= r_data[31686];
                
                r_data[31688] <= r_data[31687];
                
                r_data[31689] <= r_data[31688];
                
                r_data[31690] <= r_data[31689];
                
                r_data[31691] <= r_data[31690];
                
                r_data[31692] <= r_data[31691];
                
                r_data[31693] <= r_data[31692];
                
                r_data[31694] <= r_data[31693];
                
                r_data[31695] <= r_data[31694];
                
                r_data[31696] <= r_data[31695];
                
                r_data[31697] <= r_data[31696];
                
                r_data[31698] <= r_data[31697];
                
                r_data[31699] <= r_data[31698];
                
                r_data[31700] <= r_data[31699];
                
                r_data[31701] <= r_data[31700];
                
                r_data[31702] <= r_data[31701];
                
                r_data[31703] <= r_data[31702];
                
                r_data[31704] <= r_data[31703];
                
                r_data[31705] <= r_data[31704];
                
                r_data[31706] <= r_data[31705];
                
                r_data[31707] <= r_data[31706];
                
                r_data[31708] <= r_data[31707];
                
                r_data[31709] <= r_data[31708];
                
                r_data[31710] <= r_data[31709];
                
                r_data[31711] <= r_data[31710];
                
                r_data[31712] <= r_data[31711];
                
                r_data[31713] <= r_data[31712];
                
                r_data[31714] <= r_data[31713];
                
                r_data[31715] <= r_data[31714];
                
                r_data[31716] <= r_data[31715];
                
                r_data[31717] <= r_data[31716];
                
                r_data[31718] <= r_data[31717];
                
                r_data[31719] <= r_data[31718];
                
                r_data[31720] <= r_data[31719];
                
                r_data[31721] <= r_data[31720];
                
                r_data[31722] <= r_data[31721];
                
                r_data[31723] <= r_data[31722];
                
                r_data[31724] <= r_data[31723];
                
                r_data[31725] <= r_data[31724];
                
                r_data[31726] <= r_data[31725];
                
                r_data[31727] <= r_data[31726];
                
                r_data[31728] <= r_data[31727];
                
                r_data[31729] <= r_data[31728];
                
                r_data[31730] <= r_data[31729];
                
                r_data[31731] <= r_data[31730];
                
                r_data[31732] <= r_data[31731];
                
                r_data[31733] <= r_data[31732];
                
                r_data[31734] <= r_data[31733];
                
                r_data[31735] <= r_data[31734];
                
                r_data[31736] <= r_data[31735];
                
                r_data[31737] <= r_data[31736];
                
                r_data[31738] <= r_data[31737];
                
                r_data[31739] <= r_data[31738];
                
                r_data[31740] <= r_data[31739];
                
                r_data[31741] <= r_data[31740];
                
                r_data[31742] <= r_data[31741];
                
                r_data[31743] <= r_data[31742];
                
                r_data[31744] <= r_data[31743];
                
                r_data[31745] <= r_data[31744];
                
                r_data[31746] <= r_data[31745];
                
                r_data[31747] <= r_data[31746];
                
                r_data[31748] <= r_data[31747];
                
                r_data[31749] <= r_data[31748];
                
                r_data[31750] <= r_data[31749];
                
                r_data[31751] <= r_data[31750];
                
                r_data[31752] <= r_data[31751];
                
                r_data[31753] <= r_data[31752];
                
                r_data[31754] <= r_data[31753];
                
                r_data[31755] <= r_data[31754];
                
                r_data[31756] <= r_data[31755];
                
                r_data[31757] <= r_data[31756];
                
                r_data[31758] <= r_data[31757];
                
                r_data[31759] <= r_data[31758];
                
                r_data[31760] <= r_data[31759];
                
                r_data[31761] <= r_data[31760];
                
                r_data[31762] <= r_data[31761];
                
                r_data[31763] <= r_data[31762];
                
                r_data[31764] <= r_data[31763];
                
                r_data[31765] <= r_data[31764];
                
                r_data[31766] <= r_data[31765];
                
                r_data[31767] <= r_data[31766];
                
                r_data[31768] <= r_data[31767];
                
                r_data[31769] <= r_data[31768];
                
                r_data[31770] <= r_data[31769];
                
                r_data[31771] <= r_data[31770];
                
                r_data[31772] <= r_data[31771];
                
                r_data[31773] <= r_data[31772];
                
                r_data[31774] <= r_data[31773];
                
                r_data[31775] <= r_data[31774];
                
                r_data[31776] <= r_data[31775];
                
                r_data[31777] <= r_data[31776];
                
                r_data[31778] <= r_data[31777];
                
                r_data[31779] <= r_data[31778];
                
                r_data[31780] <= r_data[31779];
                
                r_data[31781] <= r_data[31780];
                
                r_data[31782] <= r_data[31781];
                
                r_data[31783] <= r_data[31782];
                
                r_data[31784] <= r_data[31783];
                
                r_data[31785] <= r_data[31784];
                
                r_data[31786] <= r_data[31785];
                
                r_data[31787] <= r_data[31786];
                
                r_data[31788] <= r_data[31787];
                
                r_data[31789] <= r_data[31788];
                
                r_data[31790] <= r_data[31789];
                
                r_data[31791] <= r_data[31790];
                
                r_data[31792] <= r_data[31791];
                
                r_data[31793] <= r_data[31792];
                
                r_data[31794] <= r_data[31793];
                
                r_data[31795] <= r_data[31794];
                
                r_data[31796] <= r_data[31795];
                
                r_data[31797] <= r_data[31796];
                
                r_data[31798] <= r_data[31797];
                
                r_data[31799] <= r_data[31798];
                
                r_data[31800] <= r_data[31799];
                
                r_data[31801] <= r_data[31800];
                
                r_data[31802] <= r_data[31801];
                
                r_data[31803] <= r_data[31802];
                
                r_data[31804] <= r_data[31803];
                
                r_data[31805] <= r_data[31804];
                
                r_data[31806] <= r_data[31805];
                
                r_data[31807] <= r_data[31806];
                
                r_data[31808] <= r_data[31807];
                
                r_data[31809] <= r_data[31808];
                
                r_data[31810] <= r_data[31809];
                
                r_data[31811] <= r_data[31810];
                
                r_data[31812] <= r_data[31811];
                
                r_data[31813] <= r_data[31812];
                
                r_data[31814] <= r_data[31813];
                
                r_data[31815] <= r_data[31814];
                
                r_data[31816] <= r_data[31815];
                
                r_data[31817] <= r_data[31816];
                
                r_data[31818] <= r_data[31817];
                
                r_data[31819] <= r_data[31818];
                
                r_data[31820] <= r_data[31819];
                
                r_data[31821] <= r_data[31820];
                
                r_data[31822] <= r_data[31821];
                
                r_data[31823] <= r_data[31822];
                
                r_data[31824] <= r_data[31823];
                
                r_data[31825] <= r_data[31824];
                
                r_data[31826] <= r_data[31825];
                
                r_data[31827] <= r_data[31826];
                
                r_data[31828] <= r_data[31827];
                
                r_data[31829] <= r_data[31828];
                
                r_data[31830] <= r_data[31829];
                
                r_data[31831] <= r_data[31830];
                
                r_data[31832] <= r_data[31831];
                
                r_data[31833] <= r_data[31832];
                
                r_data[31834] <= r_data[31833];
                
                r_data[31835] <= r_data[31834];
                
                r_data[31836] <= r_data[31835];
                
                r_data[31837] <= r_data[31836];
                
                r_data[31838] <= r_data[31837];
                
                r_data[31839] <= r_data[31838];
                
                r_data[31840] <= r_data[31839];
                
                r_data[31841] <= r_data[31840];
                
                r_data[31842] <= r_data[31841];
                
                r_data[31843] <= r_data[31842];
                
                r_data[31844] <= r_data[31843];
                
                r_data[31845] <= r_data[31844];
                
                r_data[31846] <= r_data[31845];
                
                r_data[31847] <= r_data[31846];
                
                r_data[31848] <= r_data[31847];
                
                r_data[31849] <= r_data[31848];
                
                r_data[31850] <= r_data[31849];
                
                r_data[31851] <= r_data[31850];
                
                r_data[31852] <= r_data[31851];
                
                r_data[31853] <= r_data[31852];
                
                r_data[31854] <= r_data[31853];
                
                r_data[31855] <= r_data[31854];
                
                r_data[31856] <= r_data[31855];
                
                r_data[31857] <= r_data[31856];
                
                r_data[31858] <= r_data[31857];
                
                r_data[31859] <= r_data[31858];
                
                r_data[31860] <= r_data[31859];
                
                r_data[31861] <= r_data[31860];
                
                r_data[31862] <= r_data[31861];
                
                r_data[31863] <= r_data[31862];
                
                r_data[31864] <= r_data[31863];
                
                r_data[31865] <= r_data[31864];
                
                r_data[31866] <= r_data[31865];
                
                r_data[31867] <= r_data[31866];
                
                r_data[31868] <= r_data[31867];
                
                r_data[31869] <= r_data[31868];
                
                r_data[31870] <= r_data[31869];
                
                r_data[31871] <= r_data[31870];
                
                r_data[31872] <= r_data[31871];
                
                r_data[31873] <= r_data[31872];
                
                r_data[31874] <= r_data[31873];
                
                r_data[31875] <= r_data[31874];
                
                r_data[31876] <= r_data[31875];
                
                r_data[31877] <= r_data[31876];
                
                r_data[31878] <= r_data[31877];
                
                r_data[31879] <= r_data[31878];
                
                r_data[31880] <= r_data[31879];
                
                r_data[31881] <= r_data[31880];
                
                r_data[31882] <= r_data[31881];
                
                r_data[31883] <= r_data[31882];
                
                r_data[31884] <= r_data[31883];
                
                r_data[31885] <= r_data[31884];
                
                r_data[31886] <= r_data[31885];
                
                r_data[31887] <= r_data[31886];
                
                r_data[31888] <= r_data[31887];
                
                r_data[31889] <= r_data[31888];
                
                r_data[31890] <= r_data[31889];
                
                r_data[31891] <= r_data[31890];
                
                r_data[31892] <= r_data[31891];
                
                r_data[31893] <= r_data[31892];
                
                r_data[31894] <= r_data[31893];
                
                r_data[31895] <= r_data[31894];
                
                r_data[31896] <= r_data[31895];
                
                r_data[31897] <= r_data[31896];
                
                r_data[31898] <= r_data[31897];
                
                r_data[31899] <= r_data[31898];
                
                r_data[31900] <= r_data[31899];
                
                r_data[31901] <= r_data[31900];
                
                r_data[31902] <= r_data[31901];
                
                r_data[31903] <= r_data[31902];
                
                r_data[31904] <= r_data[31903];
                
                r_data[31905] <= r_data[31904];
                
                r_data[31906] <= r_data[31905];
                
                r_data[31907] <= r_data[31906];
                
                r_data[31908] <= r_data[31907];
                
                r_data[31909] <= r_data[31908];
                
                r_data[31910] <= r_data[31909];
                
                r_data[31911] <= r_data[31910];
                
                r_data[31912] <= r_data[31911];
                
                r_data[31913] <= r_data[31912];
                
                r_data[31914] <= r_data[31913];
                
                r_data[31915] <= r_data[31914];
                
                r_data[31916] <= r_data[31915];
                
                r_data[31917] <= r_data[31916];
                
                r_data[31918] <= r_data[31917];
                
                r_data[31919] <= r_data[31918];
                
                r_data[31920] <= r_data[31919];
                
                r_data[31921] <= r_data[31920];
                
                r_data[31922] <= r_data[31921];
                
                r_data[31923] <= r_data[31922];
                
                r_data[31924] <= r_data[31923];
                
                r_data[31925] <= r_data[31924];
                
                r_data[31926] <= r_data[31925];
                
                r_data[31927] <= r_data[31926];
                
                r_data[31928] <= r_data[31927];
                
                r_data[31929] <= r_data[31928];
                
                r_data[31930] <= r_data[31929];
                
                r_data[31931] <= r_data[31930];
                
                r_data[31932] <= r_data[31931];
                
                r_data[31933] <= r_data[31932];
                
                r_data[31934] <= r_data[31933];
                
                r_data[31935] <= r_data[31934];
                
                r_data[31936] <= r_data[31935];
                
                r_data[31937] <= r_data[31936];
                
                r_data[31938] <= r_data[31937];
                
                r_data[31939] <= r_data[31938];
                
                r_data[31940] <= r_data[31939];
                
                r_data[31941] <= r_data[31940];
                
                r_data[31942] <= r_data[31941];
                
                r_data[31943] <= r_data[31942];
                
                r_data[31944] <= r_data[31943];
                
                r_data[31945] <= r_data[31944];
                
                r_data[31946] <= r_data[31945];
                
                r_data[31947] <= r_data[31946];
                
                r_data[31948] <= r_data[31947];
                
                r_data[31949] <= r_data[31948];
                
                r_data[31950] <= r_data[31949];
                
                r_data[31951] <= r_data[31950];
                
                r_data[31952] <= r_data[31951];
                
                r_data[31953] <= r_data[31952];
                
                r_data[31954] <= r_data[31953];
                
                r_data[31955] <= r_data[31954];
                
                r_data[31956] <= r_data[31955];
                
                r_data[31957] <= r_data[31956];
                
                r_data[31958] <= r_data[31957];
                
                r_data[31959] <= r_data[31958];
                
                r_data[31960] <= r_data[31959];
                
                r_data[31961] <= r_data[31960];
                
                r_data[31962] <= r_data[31961];
                
                r_data[31963] <= r_data[31962];
                
                r_data[31964] <= r_data[31963];
                
                r_data[31965] <= r_data[31964];
                
                r_data[31966] <= r_data[31965];
                
                r_data[31967] <= r_data[31966];
                
                r_data[31968] <= r_data[31967];
                
                r_data[31969] <= r_data[31968];
                
                r_data[31970] <= r_data[31969];
                
                r_data[31971] <= r_data[31970];
                
                r_data[31972] <= r_data[31971];
                
                r_data[31973] <= r_data[31972];
                
                r_data[31974] <= r_data[31973];
                
                r_data[31975] <= r_data[31974];
                
                r_data[31976] <= r_data[31975];
                
                r_data[31977] <= r_data[31976];
                
                r_data[31978] <= r_data[31977];
                
                r_data[31979] <= r_data[31978];
                
                r_data[31980] <= r_data[31979];
                
                r_data[31981] <= r_data[31980];
                
                r_data[31982] <= r_data[31981];
                
                r_data[31983] <= r_data[31982];
                
                r_data[31984] <= r_data[31983];
                
                r_data[31985] <= r_data[31984];
                
                r_data[31986] <= r_data[31985];
                
                r_data[31987] <= r_data[31986];
                
                r_data[31988] <= r_data[31987];
                
                r_data[31989] <= r_data[31988];
                
                r_data[31990] <= r_data[31989];
                
                r_data[31991] <= r_data[31990];
                
                r_data[31992] <= r_data[31991];
                
                r_data[31993] <= r_data[31992];
                
                r_data[31994] <= r_data[31993];
                
                r_data[31995] <= r_data[31994];
                
                r_data[31996] <= r_data[31995];
                
                r_data[31997] <= r_data[31996];
                
                r_data[31998] <= r_data[31997];
                
                r_data[31999] <= r_data[31998];
                
                r_data[32000] <= r_data[31999];
                
                r_data[32001] <= r_data[32000];
                
                r_data[32002] <= r_data[32001];
                
                r_data[32003] <= r_data[32002];
                
                r_data[32004] <= r_data[32003];
                
                r_data[32005] <= r_data[32004];
                
                r_data[32006] <= r_data[32005];
                
                r_data[32007] <= r_data[32006];
                
                r_data[32008] <= r_data[32007];
                
                r_data[32009] <= r_data[32008];
                
                r_data[32010] <= r_data[32009];
                
                r_data[32011] <= r_data[32010];
                
                r_data[32012] <= r_data[32011];
                
                r_data[32013] <= r_data[32012];
                
                r_data[32014] <= r_data[32013];
                
                r_data[32015] <= r_data[32014];
                
                r_data[32016] <= r_data[32015];
                
                r_data[32017] <= r_data[32016];
                
                r_data[32018] <= r_data[32017];
                
                r_data[32019] <= r_data[32018];
                
                r_data[32020] <= r_data[32019];
                
                r_data[32021] <= r_data[32020];
                
                r_data[32022] <= r_data[32021];
                
                r_data[32023] <= r_data[32022];
                
                r_data[32024] <= r_data[32023];
                
                r_data[32025] <= r_data[32024];
                
                r_data[32026] <= r_data[32025];
                
                r_data[32027] <= r_data[32026];
                
                r_data[32028] <= r_data[32027];
                
                r_data[32029] <= r_data[32028];
                
                r_data[32030] <= r_data[32029];
                
                r_data[32031] <= r_data[32030];
                
                r_data[32032] <= r_data[32031];
                
                r_data[32033] <= r_data[32032];
                
                r_data[32034] <= r_data[32033];
                
                r_data[32035] <= r_data[32034];
                
                r_data[32036] <= r_data[32035];
                
                r_data[32037] <= r_data[32036];
                
                r_data[32038] <= r_data[32037];
                
                r_data[32039] <= r_data[32038];
                
                r_data[32040] <= r_data[32039];
                
                r_data[32041] <= r_data[32040];
                
                r_data[32042] <= r_data[32041];
                
                r_data[32043] <= r_data[32042];
                
                r_data[32044] <= r_data[32043];
                
                r_data[32045] <= r_data[32044];
                
                r_data[32046] <= r_data[32045];
                
                r_data[32047] <= r_data[32046];
                
                r_data[32048] <= r_data[32047];
                
                r_data[32049] <= r_data[32048];
                
                r_data[32050] <= r_data[32049];
                
                r_data[32051] <= r_data[32050];
                
                r_data[32052] <= r_data[32051];
                
                r_data[32053] <= r_data[32052];
                
                r_data[32054] <= r_data[32053];
                
                r_data[32055] <= r_data[32054];
                
                r_data[32056] <= r_data[32055];
                
                r_data[32057] <= r_data[32056];
                
                r_data[32058] <= r_data[32057];
                
                r_data[32059] <= r_data[32058];
                
                r_data[32060] <= r_data[32059];
                
                r_data[32061] <= r_data[32060];
                
                r_data[32062] <= r_data[32061];
                
                r_data[32063] <= r_data[32062];
                
                r_data[32064] <= r_data[32063];
                
                r_data[32065] <= r_data[32064];
                
                r_data[32066] <= r_data[32065];
                
                r_data[32067] <= r_data[32066];
                
                r_data[32068] <= r_data[32067];
                
                r_data[32069] <= r_data[32068];
                
                r_data[32070] <= r_data[32069];
                
                r_data[32071] <= r_data[32070];
                
                r_data[32072] <= r_data[32071];
                
                r_data[32073] <= r_data[32072];
                
                r_data[32074] <= r_data[32073];
                
                r_data[32075] <= r_data[32074];
                
                r_data[32076] <= r_data[32075];
                
                r_data[32077] <= r_data[32076];
                
                r_data[32078] <= r_data[32077];
                
                r_data[32079] <= r_data[32078];
                
                r_data[32080] <= r_data[32079];
                
                r_data[32081] <= r_data[32080];
                
                r_data[32082] <= r_data[32081];
                
                r_data[32083] <= r_data[32082];
                
                r_data[32084] <= r_data[32083];
                
                r_data[32085] <= r_data[32084];
                
                r_data[32086] <= r_data[32085];
                
                r_data[32087] <= r_data[32086];
                
                r_data[32088] <= r_data[32087];
                
                r_data[32089] <= r_data[32088];
                
                r_data[32090] <= r_data[32089];
                
                r_data[32091] <= r_data[32090];
                
                r_data[32092] <= r_data[32091];
                
                r_data[32093] <= r_data[32092];
                
                r_data[32094] <= r_data[32093];
                
                r_data[32095] <= r_data[32094];
                
                r_data[32096] <= r_data[32095];
                
                r_data[32097] <= r_data[32096];
                
                r_data[32098] <= r_data[32097];
                
                r_data[32099] <= r_data[32098];
                
                r_data[32100] <= r_data[32099];
                
                r_data[32101] <= r_data[32100];
                
                r_data[32102] <= r_data[32101];
                
                r_data[32103] <= r_data[32102];
                
                r_data[32104] <= r_data[32103];
                
                r_data[32105] <= r_data[32104];
                
                r_data[32106] <= r_data[32105];
                
                r_data[32107] <= r_data[32106];
                
                r_data[32108] <= r_data[32107];
                
                r_data[32109] <= r_data[32108];
                
                r_data[32110] <= r_data[32109];
                
                r_data[32111] <= r_data[32110];
                
                r_data[32112] <= r_data[32111];
                
                r_data[32113] <= r_data[32112];
                
                r_data[32114] <= r_data[32113];
                
                r_data[32115] <= r_data[32114];
                
                r_data[32116] <= r_data[32115];
                
                r_data[32117] <= r_data[32116];
                
                r_data[32118] <= r_data[32117];
                
                r_data[32119] <= r_data[32118];
                
                r_data[32120] <= r_data[32119];
                
                r_data[32121] <= r_data[32120];
                
                r_data[32122] <= r_data[32121];
                
                r_data[32123] <= r_data[32122];
                
                r_data[32124] <= r_data[32123];
                
                r_data[32125] <= r_data[32124];
                
                r_data[32126] <= r_data[32125];
                
                r_data[32127] <= r_data[32126];
                
                r_data[32128] <= r_data[32127];
                
                r_data[32129] <= r_data[32128];
                
                r_data[32130] <= r_data[32129];
                
                r_data[32131] <= r_data[32130];
                
                r_data[32132] <= r_data[32131];
                
                r_data[32133] <= r_data[32132];
                
                r_data[32134] <= r_data[32133];
                
                r_data[32135] <= r_data[32134];
                
                r_data[32136] <= r_data[32135];
                
                r_data[32137] <= r_data[32136];
                
                r_data[32138] <= r_data[32137];
                
                r_data[32139] <= r_data[32138];
                
                r_data[32140] <= r_data[32139];
                
                r_data[32141] <= r_data[32140];
                
                r_data[32142] <= r_data[32141];
                
                r_data[32143] <= r_data[32142];
                
                r_data[32144] <= r_data[32143];
                
                r_data[32145] <= r_data[32144];
                
                r_data[32146] <= r_data[32145];
                
                r_data[32147] <= r_data[32146];
                
                r_data[32148] <= r_data[32147];
                
                r_data[32149] <= r_data[32148];
                
                r_data[32150] <= r_data[32149];
                
                r_data[32151] <= r_data[32150];
                
                r_data[32152] <= r_data[32151];
                
                r_data[32153] <= r_data[32152];
                
                r_data[32154] <= r_data[32153];
                
                r_data[32155] <= r_data[32154];
                
                r_data[32156] <= r_data[32155];
                
                r_data[32157] <= r_data[32156];
                
                r_data[32158] <= r_data[32157];
                
                r_data[32159] <= r_data[32158];
                
                r_data[32160] <= r_data[32159];
                
                r_data[32161] <= r_data[32160];
                
                r_data[32162] <= r_data[32161];
                
                r_data[32163] <= r_data[32162];
                
                r_data[32164] <= r_data[32163];
                
                r_data[32165] <= r_data[32164];
                
                r_data[32166] <= r_data[32165];
                
                r_data[32167] <= r_data[32166];
                
                r_data[32168] <= r_data[32167];
                
                r_data[32169] <= r_data[32168];
                
                r_data[32170] <= r_data[32169];
                
                r_data[32171] <= r_data[32170];
                
                r_data[32172] <= r_data[32171];
                
                r_data[32173] <= r_data[32172];
                
                r_data[32174] <= r_data[32173];
                
                r_data[32175] <= r_data[32174];
                
                r_data[32176] <= r_data[32175];
                
                r_data[32177] <= r_data[32176];
                
                r_data[32178] <= r_data[32177];
                
                r_data[32179] <= r_data[32178];
                
                r_data[32180] <= r_data[32179];
                
                r_data[32181] <= r_data[32180];
                
                r_data[32182] <= r_data[32181];
                
                r_data[32183] <= r_data[32182];
                
                r_data[32184] <= r_data[32183];
                
                r_data[32185] <= r_data[32184];
                
                r_data[32186] <= r_data[32185];
                
                r_data[32187] <= r_data[32186];
                
                r_data[32188] <= r_data[32187];
                
                r_data[32189] <= r_data[32188];
                
                r_data[32190] <= r_data[32189];
                
                r_data[32191] <= r_data[32190];
                
                r_data[32192] <= r_data[32191];
                
                r_data[32193] <= r_data[32192];
                
                r_data[32194] <= r_data[32193];
                
                r_data[32195] <= r_data[32194];
                
                r_data[32196] <= r_data[32195];
                
                r_data[32197] <= r_data[32196];
                
                r_data[32198] <= r_data[32197];
                
                r_data[32199] <= r_data[32198];
                
                r_data[32200] <= r_data[32199];
                
                r_data[32201] <= r_data[32200];
                
                r_data[32202] <= r_data[32201];
                
                r_data[32203] <= r_data[32202];
                
                r_data[32204] <= r_data[32203];
                
                r_data[32205] <= r_data[32204];
                
                r_data[32206] <= r_data[32205];
                
                r_data[32207] <= r_data[32206];
                
                r_data[32208] <= r_data[32207];
                
                r_data[32209] <= r_data[32208];
                
                r_data[32210] <= r_data[32209];
                
                r_data[32211] <= r_data[32210];
                
                r_data[32212] <= r_data[32211];
                
                r_data[32213] <= r_data[32212];
                
                r_data[32214] <= r_data[32213];
                
                r_data[32215] <= r_data[32214];
                
                r_data[32216] <= r_data[32215];
                
                r_data[32217] <= r_data[32216];
                
                r_data[32218] <= r_data[32217];
                
                r_data[32219] <= r_data[32218];
                
                r_data[32220] <= r_data[32219];
                
                r_data[32221] <= r_data[32220];
                
                r_data[32222] <= r_data[32221];
                
                r_data[32223] <= r_data[32222];
                
                r_data[32224] <= r_data[32223];
                
                r_data[32225] <= r_data[32224];
                
                r_data[32226] <= r_data[32225];
                
                r_data[32227] <= r_data[32226];
                
                r_data[32228] <= r_data[32227];
                
                r_data[32229] <= r_data[32228];
                
                r_data[32230] <= r_data[32229];
                
                r_data[32231] <= r_data[32230];
                
                r_data[32232] <= r_data[32231];
                
                r_data[32233] <= r_data[32232];
                
                r_data[32234] <= r_data[32233];
                
                r_data[32235] <= r_data[32234];
                
                r_data[32236] <= r_data[32235];
                
                r_data[32237] <= r_data[32236];
                
                r_data[32238] <= r_data[32237];
                
                r_data[32239] <= r_data[32238];
                
                r_data[32240] <= r_data[32239];
                
                r_data[32241] <= r_data[32240];
                
                r_data[32242] <= r_data[32241];
                
                r_data[32243] <= r_data[32242];
                
                r_data[32244] <= r_data[32243];
                
                r_data[32245] <= r_data[32244];
                
                r_data[32246] <= r_data[32245];
                
                r_data[32247] <= r_data[32246];
                
                r_data[32248] <= r_data[32247];
                
                r_data[32249] <= r_data[32248];
                
                r_data[32250] <= r_data[32249];
                
                r_data[32251] <= r_data[32250];
                
                r_data[32252] <= r_data[32251];
                
                r_data[32253] <= r_data[32252];
                
                r_data[32254] <= r_data[32253];
                
                r_data[32255] <= r_data[32254];
                
                r_data[32256] <= r_data[32255];
                
                r_data[32257] <= r_data[32256];
                
                r_data[32258] <= r_data[32257];
                
                r_data[32259] <= r_data[32258];
                
                r_data[32260] <= r_data[32259];
                
                r_data[32261] <= r_data[32260];
                
                r_data[32262] <= r_data[32261];
                
                r_data[32263] <= r_data[32262];
                
                r_data[32264] <= r_data[32263];
                
                r_data[32265] <= r_data[32264];
                
                r_data[32266] <= r_data[32265];
                
                r_data[32267] <= r_data[32266];
                
                r_data[32268] <= r_data[32267];
                
                r_data[32269] <= r_data[32268];
                
                r_data[32270] <= r_data[32269];
                
                r_data[32271] <= r_data[32270];
                
                r_data[32272] <= r_data[32271];
                
                r_data[32273] <= r_data[32272];
                
                r_data[32274] <= r_data[32273];
                
                r_data[32275] <= r_data[32274];
                
                r_data[32276] <= r_data[32275];
                
                r_data[32277] <= r_data[32276];
                
                r_data[32278] <= r_data[32277];
                
                r_data[32279] <= r_data[32278];
                
                r_data[32280] <= r_data[32279];
                
                r_data[32281] <= r_data[32280];
                
                r_data[32282] <= r_data[32281];
                
                r_data[32283] <= r_data[32282];
                
                r_data[32284] <= r_data[32283];
                
                r_data[32285] <= r_data[32284];
                
                r_data[32286] <= r_data[32285];
                
                r_data[32287] <= r_data[32286];
                
                r_data[32288] <= r_data[32287];
                
                r_data[32289] <= r_data[32288];
                
                r_data[32290] <= r_data[32289];
                
                r_data[32291] <= r_data[32290];
                
                r_data[32292] <= r_data[32291];
                
                r_data[32293] <= r_data[32292];
                
                r_data[32294] <= r_data[32293];
                
                r_data[32295] <= r_data[32294];
                
                r_data[32296] <= r_data[32295];
                
                r_data[32297] <= r_data[32296];
                
                r_data[32298] <= r_data[32297];
                
                r_data[32299] <= r_data[32298];
                
                r_data[32300] <= r_data[32299];
                
                r_data[32301] <= r_data[32300];
                
                r_data[32302] <= r_data[32301];
                
                r_data[32303] <= r_data[32302];
                
                r_data[32304] <= r_data[32303];
                
                r_data[32305] <= r_data[32304];
                
                r_data[32306] <= r_data[32305];
                
                r_data[32307] <= r_data[32306];
                
                r_data[32308] <= r_data[32307];
                
                r_data[32309] <= r_data[32308];
                
                r_data[32310] <= r_data[32309];
                
                r_data[32311] <= r_data[32310];
                
                r_data[32312] <= r_data[32311];
                
                r_data[32313] <= r_data[32312];
                
                r_data[32314] <= r_data[32313];
                
                r_data[32315] <= r_data[32314];
                
                r_data[32316] <= r_data[32315];
                
                r_data[32317] <= r_data[32316];
                
                r_data[32318] <= r_data[32317];
                
                r_data[32319] <= r_data[32318];
                
                r_data[32320] <= r_data[32319];
                
                r_data[32321] <= r_data[32320];
                
                r_data[32322] <= r_data[32321];
                
                r_data[32323] <= r_data[32322];
                
                r_data[32324] <= r_data[32323];
                
                r_data[32325] <= r_data[32324];
                
                r_data[32326] <= r_data[32325];
                
                r_data[32327] <= r_data[32326];
                
                r_data[32328] <= r_data[32327];
                
                r_data[32329] <= r_data[32328];
                
                r_data[32330] <= r_data[32329];
                
                r_data[32331] <= r_data[32330];
                
                r_data[32332] <= r_data[32331];
                
                r_data[32333] <= r_data[32332];
                
                r_data[32334] <= r_data[32333];
                
                r_data[32335] <= r_data[32334];
                
                r_data[32336] <= r_data[32335];
                
                r_data[32337] <= r_data[32336];
                
                r_data[32338] <= r_data[32337];
                
                r_data[32339] <= r_data[32338];
                
                r_data[32340] <= r_data[32339];
                
                r_data[32341] <= r_data[32340];
                
                r_data[32342] <= r_data[32341];
                
                r_data[32343] <= r_data[32342];
                
                r_data[32344] <= r_data[32343];
                
                r_data[32345] <= r_data[32344];
                
                r_data[32346] <= r_data[32345];
                
                r_data[32347] <= r_data[32346];
                
                r_data[32348] <= r_data[32347];
                
                r_data[32349] <= r_data[32348];
                
                r_data[32350] <= r_data[32349];
                
                r_data[32351] <= r_data[32350];
                
                r_data[32352] <= r_data[32351];
                
                r_data[32353] <= r_data[32352];
                
                r_data[32354] <= r_data[32353];
                
                r_data[32355] <= r_data[32354];
                
                r_data[32356] <= r_data[32355];
                
                r_data[32357] <= r_data[32356];
                
                r_data[32358] <= r_data[32357];
                
                r_data[32359] <= r_data[32358];
                
                r_data[32360] <= r_data[32359];
                
                r_data[32361] <= r_data[32360];
                
                r_data[32362] <= r_data[32361];
                
                r_data[32363] <= r_data[32362];
                
                r_data[32364] <= r_data[32363];
                
                r_data[32365] <= r_data[32364];
                
                r_data[32366] <= r_data[32365];
                
                r_data[32367] <= r_data[32366];
                
                r_data[32368] <= r_data[32367];
                
                r_data[32369] <= r_data[32368];
                
                r_data[32370] <= r_data[32369];
                
                r_data[32371] <= r_data[32370];
                
                r_data[32372] <= r_data[32371];
                
                r_data[32373] <= r_data[32372];
                
                r_data[32374] <= r_data[32373];
                
                r_data[32375] <= r_data[32374];
                
                r_data[32376] <= r_data[32375];
                
                r_data[32377] <= r_data[32376];
                
                r_data[32378] <= r_data[32377];
                
                r_data[32379] <= r_data[32378];
                
                r_data[32380] <= r_data[32379];
                
                r_data[32381] <= r_data[32380];
                
                r_data[32382] <= r_data[32381];
                
                r_data[32383] <= r_data[32382];
                
                r_data[32384] <= r_data[32383];
                
                r_data[32385] <= r_data[32384];
                
                r_data[32386] <= r_data[32385];
                
                r_data[32387] <= r_data[32386];
                
                r_data[32388] <= r_data[32387];
                
                r_data[32389] <= r_data[32388];
                
                r_data[32390] <= r_data[32389];
                
                r_data[32391] <= r_data[32390];
                
                r_data[32392] <= r_data[32391];
                
                r_data[32393] <= r_data[32392];
                
                r_data[32394] <= r_data[32393];
                
                r_data[32395] <= r_data[32394];
                
                r_data[32396] <= r_data[32395];
                
                r_data[32397] <= r_data[32396];
                
                r_data[32398] <= r_data[32397];
                
                r_data[32399] <= r_data[32398];
                
                r_data[32400] <= r_data[32399];
                
                r_data[32401] <= r_data[32400];
                
                r_data[32402] <= r_data[32401];
                
                r_data[32403] <= r_data[32402];
                
                r_data[32404] <= r_data[32403];
                
                r_data[32405] <= r_data[32404];
                
                r_data[32406] <= r_data[32405];
                
                r_data[32407] <= r_data[32406];
                
                r_data[32408] <= r_data[32407];
                
                r_data[32409] <= r_data[32408];
                
                r_data[32410] <= r_data[32409];
                
                r_data[32411] <= r_data[32410];
                
                r_data[32412] <= r_data[32411];
                
                r_data[32413] <= r_data[32412];
                
                r_data[32414] <= r_data[32413];
                
                r_data[32415] <= r_data[32414];
                
                r_data[32416] <= r_data[32415];
                
                r_data[32417] <= r_data[32416];
                
                r_data[32418] <= r_data[32417];
                
                r_data[32419] <= r_data[32418];
                
                r_data[32420] <= r_data[32419];
                
                r_data[32421] <= r_data[32420];
                
                r_data[32422] <= r_data[32421];
                
                r_data[32423] <= r_data[32422];
                
                r_data[32424] <= r_data[32423];
                
                r_data[32425] <= r_data[32424];
                
                r_data[32426] <= r_data[32425];
                
                r_data[32427] <= r_data[32426];
                
                r_data[32428] <= r_data[32427];
                
                r_data[32429] <= r_data[32428];
                
                r_data[32430] <= r_data[32429];
                
                r_data[32431] <= r_data[32430];
                
                r_data[32432] <= r_data[32431];
                
                r_data[32433] <= r_data[32432];
                
                r_data[32434] <= r_data[32433];
                
                r_data[32435] <= r_data[32434];
                
                r_data[32436] <= r_data[32435];
                
                r_data[32437] <= r_data[32436];
                
                r_data[32438] <= r_data[32437];
                
                r_data[32439] <= r_data[32438];
                
                r_data[32440] <= r_data[32439];
                
                r_data[32441] <= r_data[32440];
                
                r_data[32442] <= r_data[32441];
                
                r_data[32443] <= r_data[32442];
                
                r_data[32444] <= r_data[32443];
                
                r_data[32445] <= r_data[32444];
                
                r_data[32446] <= r_data[32445];
                
                r_data[32447] <= r_data[32446];
                
                r_data[32448] <= r_data[32447];
                
                r_data[32449] <= r_data[32448];
                
                r_data[32450] <= r_data[32449];
                
                r_data[32451] <= r_data[32450];
                
                r_data[32452] <= r_data[32451];
                
                r_data[32453] <= r_data[32452];
                
                r_data[32454] <= r_data[32453];
                
                r_data[32455] <= r_data[32454];
                
                r_data[32456] <= r_data[32455];
                
                r_data[32457] <= r_data[32456];
                
                r_data[32458] <= r_data[32457];
                
                r_data[32459] <= r_data[32458];
                
                r_data[32460] <= r_data[32459];
                
                r_data[32461] <= r_data[32460];
                
                r_data[32462] <= r_data[32461];
                
                r_data[32463] <= r_data[32462];
                
                r_data[32464] <= r_data[32463];
                
                r_data[32465] <= r_data[32464];
                
                r_data[32466] <= r_data[32465];
                
                r_data[32467] <= r_data[32466];
                
                r_data[32468] <= r_data[32467];
                
                r_data[32469] <= r_data[32468];
                
                r_data[32470] <= r_data[32469];
                
                r_data[32471] <= r_data[32470];
                
                r_data[32472] <= r_data[32471];
                
                r_data[32473] <= r_data[32472];
                
                r_data[32474] <= r_data[32473];
                
                r_data[32475] <= r_data[32474];
                
                r_data[32476] <= r_data[32475];
                
                r_data[32477] <= r_data[32476];
                
                r_data[32478] <= r_data[32477];
                
                r_data[32479] <= r_data[32478];
                
                r_data[32480] <= r_data[32479];
                
                r_data[32481] <= r_data[32480];
                
                r_data[32482] <= r_data[32481];
                
                r_data[32483] <= r_data[32482];
                
                r_data[32484] <= r_data[32483];
                
                r_data[32485] <= r_data[32484];
                
                r_data[32486] <= r_data[32485];
                
                r_data[32487] <= r_data[32486];
                
                r_data[32488] <= r_data[32487];
                
                r_data[32489] <= r_data[32488];
                
                r_data[32490] <= r_data[32489];
                
                r_data[32491] <= r_data[32490];
                
                r_data[32492] <= r_data[32491];
                
                r_data[32493] <= r_data[32492];
                
                r_data[32494] <= r_data[32493];
                
                r_data[32495] <= r_data[32494];
                
                r_data[32496] <= r_data[32495];
                
                r_data[32497] <= r_data[32496];
                
                r_data[32498] <= r_data[32497];
                
                r_data[32499] <= r_data[32498];
                
                r_data[32500] <= r_data[32499];
                
                r_data[32501] <= r_data[32500];
                
                r_data[32502] <= r_data[32501];
                
                r_data[32503] <= r_data[32502];
                
                r_data[32504] <= r_data[32503];
                
                r_data[32505] <= r_data[32504];
                
                r_data[32506] <= r_data[32505];
                
                r_data[32507] <= r_data[32506];
                
                r_data[32508] <= r_data[32507];
                
                r_data[32509] <= r_data[32508];
                
                r_data[32510] <= r_data[32509];
                
                r_data[32511] <= r_data[32510];
                
                r_data[32512] <= r_data[32511];
                
                r_data[32513] <= r_data[32512];
                
                r_data[32514] <= r_data[32513];
                
                r_data[32515] <= r_data[32514];
                
                r_data[32516] <= r_data[32515];
                
                r_data[32517] <= r_data[32516];
                
                r_data[32518] <= r_data[32517];
                
                r_data[32519] <= r_data[32518];
                
                r_data[32520] <= r_data[32519];
                
                r_data[32521] <= r_data[32520];
                
                r_data[32522] <= r_data[32521];
                
                r_data[32523] <= r_data[32522];
                
                r_data[32524] <= r_data[32523];
                
                r_data[32525] <= r_data[32524];
                
                r_data[32526] <= r_data[32525];
                
                r_data[32527] <= r_data[32526];
                
                r_data[32528] <= r_data[32527];
                
                r_data[32529] <= r_data[32528];
                
                r_data[32530] <= r_data[32529];
                
                r_data[32531] <= r_data[32530];
                
                r_data[32532] <= r_data[32531];
                
                r_data[32533] <= r_data[32532];
                
                r_data[32534] <= r_data[32533];
                
                r_data[32535] <= r_data[32534];
                
                r_data[32536] <= r_data[32535];
                
                r_data[32537] <= r_data[32536];
                
                r_data[32538] <= r_data[32537];
                
                r_data[32539] <= r_data[32538];
                
                r_data[32540] <= r_data[32539];
                
                r_data[32541] <= r_data[32540];
                
                r_data[32542] <= r_data[32541];
                
                r_data[32543] <= r_data[32542];
                
                r_data[32544] <= r_data[32543];
                
                r_data[32545] <= r_data[32544];
                
                r_data[32546] <= r_data[32545];
                
                r_data[32547] <= r_data[32546];
                
                r_data[32548] <= r_data[32547];
                
                r_data[32549] <= r_data[32548];
                
                r_data[32550] <= r_data[32549];
                
                r_data[32551] <= r_data[32550];
                
                r_data[32552] <= r_data[32551];
                
                r_data[32553] <= r_data[32552];
                
                r_data[32554] <= r_data[32553];
                
                r_data[32555] <= r_data[32554];
                
                r_data[32556] <= r_data[32555];
                
                r_data[32557] <= r_data[32556];
                
                r_data[32558] <= r_data[32557];
                
                r_data[32559] <= r_data[32558];
                
                r_data[32560] <= r_data[32559];
                
                r_data[32561] <= r_data[32560];
                
                r_data[32562] <= r_data[32561];
                
                r_data[32563] <= r_data[32562];
                
                r_data[32564] <= r_data[32563];
                
                r_data[32565] <= r_data[32564];
                
                r_data[32566] <= r_data[32565];
                
                r_data[32567] <= r_data[32566];
                
                r_data[32568] <= r_data[32567];
                
                r_data[32569] <= r_data[32568];
                
                r_data[32570] <= r_data[32569];
                
                r_data[32571] <= r_data[32570];
                
                r_data[32572] <= r_data[32571];
                
                r_data[32573] <= r_data[32572];
                
                r_data[32574] <= r_data[32573];
                
                r_data[32575] <= r_data[32574];
                
                r_data[32576] <= r_data[32575];
                
                r_data[32577] <= r_data[32576];
                
                r_data[32578] <= r_data[32577];
                
                r_data[32579] <= r_data[32578];
                
                r_data[32580] <= r_data[32579];
                
                r_data[32581] <= r_data[32580];
                
                r_data[32582] <= r_data[32581];
                
                r_data[32583] <= r_data[32582];
                
                r_data[32584] <= r_data[32583];
                
                r_data[32585] <= r_data[32584];
                
                r_data[32586] <= r_data[32585];
                
                r_data[32587] <= r_data[32586];
                
                r_data[32588] <= r_data[32587];
                
                r_data[32589] <= r_data[32588];
                
                r_data[32590] <= r_data[32589];
                
                r_data[32591] <= r_data[32590];
                
                r_data[32592] <= r_data[32591];
                
                r_data[32593] <= r_data[32592];
                
                r_data[32594] <= r_data[32593];
                
                r_data[32595] <= r_data[32594];
                
                r_data[32596] <= r_data[32595];
                
                r_data[32597] <= r_data[32596];
                
                r_data[32598] <= r_data[32597];
                
                r_data[32599] <= r_data[32598];
                
                r_data[32600] <= r_data[32599];
                
                r_data[32601] <= r_data[32600];
                
                r_data[32602] <= r_data[32601];
                
                r_data[32603] <= r_data[32602];
                
                r_data[32604] <= r_data[32603];
                
                r_data[32605] <= r_data[32604];
                
                r_data[32606] <= r_data[32605];
                
                r_data[32607] <= r_data[32606];
                
                r_data[32608] <= r_data[32607];
                
                r_data[32609] <= r_data[32608];
                
                r_data[32610] <= r_data[32609];
                
                r_data[32611] <= r_data[32610];
                
                r_data[32612] <= r_data[32611];
                
                r_data[32613] <= r_data[32612];
                
                r_data[32614] <= r_data[32613];
                
                r_data[32615] <= r_data[32614];
                
                r_data[32616] <= r_data[32615];
                
                r_data[32617] <= r_data[32616];
                
                r_data[32618] <= r_data[32617];
                
                r_data[32619] <= r_data[32618];
                
                r_data[32620] <= r_data[32619];
                
                r_data[32621] <= r_data[32620];
                
                r_data[32622] <= r_data[32621];
                
                r_data[32623] <= r_data[32622];
                
                r_data[32624] <= r_data[32623];
                
                r_data[32625] <= r_data[32624];
                
                r_data[32626] <= r_data[32625];
                
                r_data[32627] <= r_data[32626];
                
                r_data[32628] <= r_data[32627];
                
                r_data[32629] <= r_data[32628];
                
                r_data[32630] <= r_data[32629];
                
                r_data[32631] <= r_data[32630];
                
                r_data[32632] <= r_data[32631];
                
                r_data[32633] <= r_data[32632];
                
                r_data[32634] <= r_data[32633];
                
                r_data[32635] <= r_data[32634];
                
                r_data[32636] <= r_data[32635];
                
                r_data[32637] <= r_data[32636];
                
                r_data[32638] <= r_data[32637];
                
                r_data[32639] <= r_data[32638];
                
                r_data[32640] <= r_data[32639];
                
                r_data[32641] <= r_data[32640];
                
                r_data[32642] <= r_data[32641];
                
                r_data[32643] <= r_data[32642];
                
                r_data[32644] <= r_data[32643];
                
                r_data[32645] <= r_data[32644];
                
                r_data[32646] <= r_data[32645];
                
                r_data[32647] <= r_data[32646];
                
                r_data[32648] <= r_data[32647];
                
                r_data[32649] <= r_data[32648];
                
                r_data[32650] <= r_data[32649];
                
                r_data[32651] <= r_data[32650];
                
                r_data[32652] <= r_data[32651];
                
                r_data[32653] <= r_data[32652];
                
                r_data[32654] <= r_data[32653];
                
                r_data[32655] <= r_data[32654];
                
                r_data[32656] <= r_data[32655];
                
                r_data[32657] <= r_data[32656];
                
                r_data[32658] <= r_data[32657];
                
                r_data[32659] <= r_data[32658];
                
                r_data[32660] <= r_data[32659];
                
                r_data[32661] <= r_data[32660];
                
                r_data[32662] <= r_data[32661];
                
                r_data[32663] <= r_data[32662];
                
                r_data[32664] <= r_data[32663];
                
                r_data[32665] <= r_data[32664];
                
                r_data[32666] <= r_data[32665];
                
                r_data[32667] <= r_data[32666];
                
                r_data[32668] <= r_data[32667];
                
                r_data[32669] <= r_data[32668];
                
                r_data[32670] <= r_data[32669];
                
                r_data[32671] <= r_data[32670];
                
                r_data[32672] <= r_data[32671];
                
                r_data[32673] <= r_data[32672];
                
                r_data[32674] <= r_data[32673];
                
                r_data[32675] <= r_data[32674];
                
                r_data[32676] <= r_data[32675];
                
                r_data[32677] <= r_data[32676];
                
                r_data[32678] <= r_data[32677];
                
                r_data[32679] <= r_data[32678];
                
                r_data[32680] <= r_data[32679];
                
                r_data[32681] <= r_data[32680];
                
                r_data[32682] <= r_data[32681];
                
                r_data[32683] <= r_data[32682];
                
                r_data[32684] <= r_data[32683];
                
                r_data[32685] <= r_data[32684];
                
                r_data[32686] <= r_data[32685];
                
                r_data[32687] <= r_data[32686];
                
                r_data[32688] <= r_data[32687];
                
                r_data[32689] <= r_data[32688];
                
                r_data[32690] <= r_data[32689];
                
                r_data[32691] <= r_data[32690];
                
                r_data[32692] <= r_data[32691];
                
                r_data[32693] <= r_data[32692];
                
                r_data[32694] <= r_data[32693];
                
                r_data[32695] <= r_data[32694];
                
                r_data[32696] <= r_data[32695];
                
                r_data[32697] <= r_data[32696];
                
                r_data[32698] <= r_data[32697];
                
                r_data[32699] <= r_data[32698];
                
                r_data[32700] <= r_data[32699];
                
                r_data[32701] <= r_data[32700];
                
                r_data[32702] <= r_data[32701];
                
                r_data[32703] <= r_data[32702];
                
                r_data[32704] <= r_data[32703];
                
                r_data[32705] <= r_data[32704];
                
                r_data[32706] <= r_data[32705];
                
                r_data[32707] <= r_data[32706];
                
                r_data[32708] <= r_data[32707];
                
                r_data[32709] <= r_data[32708];
                
                r_data[32710] <= r_data[32709];
                
                r_data[32711] <= r_data[32710];
                
                r_data[32712] <= r_data[32711];
                
                r_data[32713] <= r_data[32712];
                
                r_data[32714] <= r_data[32713];
                
                r_data[32715] <= r_data[32714];
                
                r_data[32716] <= r_data[32715];
                
                r_data[32717] <= r_data[32716];
                
                r_data[32718] <= r_data[32717];
                
                r_data[32719] <= r_data[32718];
                
                r_data[32720] <= r_data[32719];
                
                r_data[32721] <= r_data[32720];
                
                r_data[32722] <= r_data[32721];
                
                r_data[32723] <= r_data[32722];
                
                r_data[32724] <= r_data[32723];
                
                r_data[32725] <= r_data[32724];
                
                r_data[32726] <= r_data[32725];
                
                r_data[32727] <= r_data[32726];
                
                r_data[32728] <= r_data[32727];
                
                r_data[32729] <= r_data[32728];
                
                r_data[32730] <= r_data[32729];
                
                r_data[32731] <= r_data[32730];
                
                r_data[32732] <= r_data[32731];
                
                r_data[32733] <= r_data[32732];
                
                r_data[32734] <= r_data[32733];
                
                r_data[32735] <= r_data[32734];
                
                r_data[32736] <= r_data[32735];
                
                r_data[32737] <= r_data[32736];
                
                r_data[32738] <= r_data[32737];
                
                r_data[32739] <= r_data[32738];
                
                r_data[32740] <= r_data[32739];
                
                r_data[32741] <= r_data[32740];
                
                r_data[32742] <= r_data[32741];
                
                r_data[32743] <= r_data[32742];
                
                r_data[32744] <= r_data[32743];
                
                r_data[32745] <= r_data[32744];
                
                r_data[32746] <= r_data[32745];
                
                r_data[32747] <= r_data[32746];
                
                r_data[32748] <= r_data[32747];
                
                r_data[32749] <= r_data[32748];
                
                r_data[32750] <= r_data[32749];
                
                r_data[32751] <= r_data[32750];
                
                r_data[32752] <= r_data[32751];
                
                r_data[32753] <= r_data[32752];
                
                r_data[32754] <= r_data[32753];
                
                r_data[32755] <= r_data[32754];
                
                r_data[32756] <= r_data[32755];
                
                r_data[32757] <= r_data[32756];
                
                r_data[32758] <= r_data[32757];
                
                r_data[32759] <= r_data[32758];
                
                r_data[32760] <= r_data[32759];
                
                r_data[32761] <= r_data[32760];
                
                r_data[32762] <= r_data[32761];
                
                r_data[32763] <= r_data[32762];
                
                r_data[32764] <= r_data[32763];
                
                r_data[32765] <= r_data[32764];
                
                r_data[32766] <= r_data[32765];
                
                r_data[32767] <= r_data[32766];
                
                r_data[32768] <= r_data[32767];
                
                r_data[32769] <= r_data[32768];
                
                r_data[32770] <= r_data[32769];
                
                r_data[32771] <= r_data[32770];
                
                r_data[32772] <= r_data[32771];
                
                r_data[32773] <= r_data[32772];
                
                r_data[32774] <= r_data[32773];
                
                r_data[32775] <= r_data[32774];
                
                r_data[32776] <= r_data[32775];
                
                r_data[32777] <= r_data[32776];
                
                r_data[32778] <= r_data[32777];
                
                r_data[32779] <= r_data[32778];
                
                r_data[32780] <= r_data[32779];
                
                r_data[32781] <= r_data[32780];
                
                r_data[32782] <= r_data[32781];
                
                r_data[32783] <= r_data[32782];
                
                r_data[32784] <= r_data[32783];
                
                r_data[32785] <= r_data[32784];
                
                r_data[32786] <= r_data[32785];
                
                r_data[32787] <= r_data[32786];
                
                r_data[32788] <= r_data[32787];
                
                r_data[32789] <= r_data[32788];
                
                r_data[32790] <= r_data[32789];
                
                r_data[32791] <= r_data[32790];
                
                r_data[32792] <= r_data[32791];
                
                r_data[32793] <= r_data[32792];
                
                r_data[32794] <= r_data[32793];
                
                r_data[32795] <= r_data[32794];
                
                r_data[32796] <= r_data[32795];
                
                r_data[32797] <= r_data[32796];
                
                r_data[32798] <= r_data[32797];
                
                r_data[32799] <= r_data[32798];
                
                r_data[32800] <= r_data[32799];
                
                r_data[32801] <= r_data[32800];
                
                r_data[32802] <= r_data[32801];
                
                r_data[32803] <= r_data[32802];
                
                r_data[32804] <= r_data[32803];
                
                r_data[32805] <= r_data[32804];
                
                r_data[32806] <= r_data[32805];
                
                r_data[32807] <= r_data[32806];
                
                r_data[32808] <= r_data[32807];
                
                r_data[32809] <= r_data[32808];
                
                r_data[32810] <= r_data[32809];
                
                r_data[32811] <= r_data[32810];
                
                r_data[32812] <= r_data[32811];
                
                r_data[32813] <= r_data[32812];
                
                r_data[32814] <= r_data[32813];
                
                r_data[32815] <= r_data[32814];
                
                r_data[32816] <= r_data[32815];
                
                r_data[32817] <= r_data[32816];
                
                r_data[32818] <= r_data[32817];
                
                r_data[32819] <= r_data[32818];
                
                r_data[32820] <= r_data[32819];
                
                r_data[32821] <= r_data[32820];
                
                r_data[32822] <= r_data[32821];
                
                r_data[32823] <= r_data[32822];
                
                r_data[32824] <= r_data[32823];
                
                r_data[32825] <= r_data[32824];
                
                r_data[32826] <= r_data[32825];
                
                r_data[32827] <= r_data[32826];
                
                r_data[32828] <= r_data[32827];
                
                r_data[32829] <= r_data[32828];
                
                r_data[32830] <= r_data[32829];
                
                r_data[32831] <= r_data[32830];
                
                r_data[32832] <= r_data[32831];
                
                r_data[32833] <= r_data[32832];
                
                r_data[32834] <= r_data[32833];
                
                r_data[32835] <= r_data[32834];
                
                r_data[32836] <= r_data[32835];
                
                r_data[32837] <= r_data[32836];
                
                r_data[32838] <= r_data[32837];
                
                r_data[32839] <= r_data[32838];
                
                r_data[32840] <= r_data[32839];
                
                r_data[32841] <= r_data[32840];
                
                r_data[32842] <= r_data[32841];
                
                r_data[32843] <= r_data[32842];
                
                r_data[32844] <= r_data[32843];
                
                r_data[32845] <= r_data[32844];
                
                r_data[32846] <= r_data[32845];
                
                r_data[32847] <= r_data[32846];
                
                r_data[32848] <= r_data[32847];
                
                r_data[32849] <= r_data[32848];
                
                r_data[32850] <= r_data[32849];
                
                r_data[32851] <= r_data[32850];
                
                r_data[32852] <= r_data[32851];
                
                r_data[32853] <= r_data[32852];
                
                r_data[32854] <= r_data[32853];
                
                r_data[32855] <= r_data[32854];
                
                r_data[32856] <= r_data[32855];
                
                r_data[32857] <= r_data[32856];
                
                r_data[32858] <= r_data[32857];
                
                r_data[32859] <= r_data[32858];
                
                r_data[32860] <= r_data[32859];
                
                r_data[32861] <= r_data[32860];
                
                r_data[32862] <= r_data[32861];
                
                r_data[32863] <= r_data[32862];
                
                r_data[32864] <= r_data[32863];
                
                r_data[32865] <= r_data[32864];
                
                r_data[32866] <= r_data[32865];
                
                r_data[32867] <= r_data[32866];
                
                r_data[32868] <= r_data[32867];
                
                r_data[32869] <= r_data[32868];
                
                r_data[32870] <= r_data[32869];
                
                r_data[32871] <= r_data[32870];
                
                r_data[32872] <= r_data[32871];
                
                r_data[32873] <= r_data[32872];
                
                r_data[32874] <= r_data[32873];
                
                r_data[32875] <= r_data[32874];
                
                r_data[32876] <= r_data[32875];
                
                r_data[32877] <= r_data[32876];
                
                r_data[32878] <= r_data[32877];
                
                r_data[32879] <= r_data[32878];
                
                r_data[32880] <= r_data[32879];
                
                r_data[32881] <= r_data[32880];
                
                r_data[32882] <= r_data[32881];
                
                r_data[32883] <= r_data[32882];
                
                r_data[32884] <= r_data[32883];
                
                r_data[32885] <= r_data[32884];
                
                r_data[32886] <= r_data[32885];
                
                r_data[32887] <= r_data[32886];
                
                r_data[32888] <= r_data[32887];
                
                r_data[32889] <= r_data[32888];
                
                r_data[32890] <= r_data[32889];
                
                r_data[32891] <= r_data[32890];
                
                r_data[32892] <= r_data[32891];
                
                r_data[32893] <= r_data[32892];
                
                r_data[32894] <= r_data[32893];
                
                r_data[32895] <= r_data[32894];
                
                r_data[32896] <= r_data[32895];
                
                r_data[32897] <= r_data[32896];
                
                r_data[32898] <= r_data[32897];
                
                r_data[32899] <= r_data[32898];
                
                r_data[32900] <= r_data[32899];
                
                r_data[32901] <= r_data[32900];
                
                r_data[32902] <= r_data[32901];
                
                r_data[32903] <= r_data[32902];
                
                r_data[32904] <= r_data[32903];
                
                r_data[32905] <= r_data[32904];
                
                r_data[32906] <= r_data[32905];
                
                r_data[32907] <= r_data[32906];
                
                r_data[32908] <= r_data[32907];
                
                r_data[32909] <= r_data[32908];
                
                r_data[32910] <= r_data[32909];
                
                r_data[32911] <= r_data[32910];
                
                r_data[32912] <= r_data[32911];
                
                r_data[32913] <= r_data[32912];
                
                r_data[32914] <= r_data[32913];
                
                r_data[32915] <= r_data[32914];
                
                r_data[32916] <= r_data[32915];
                
                r_data[32917] <= r_data[32916];
                
                r_data[32918] <= r_data[32917];
                
                r_data[32919] <= r_data[32918];
                
                r_data[32920] <= r_data[32919];
                
                r_data[32921] <= r_data[32920];
                
                r_data[32922] <= r_data[32921];
                
                r_data[32923] <= r_data[32922];
                
                r_data[32924] <= r_data[32923];
                
                r_data[32925] <= r_data[32924];
                
                r_data[32926] <= r_data[32925];
                
                r_data[32927] <= r_data[32926];
                
                r_data[32928] <= r_data[32927];
                
                r_data[32929] <= r_data[32928];
                
                r_data[32930] <= r_data[32929];
                
                r_data[32931] <= r_data[32930];
                
                r_data[32932] <= r_data[32931];
                
                r_data[32933] <= r_data[32932];
                
                r_data[32934] <= r_data[32933];
                
                r_data[32935] <= r_data[32934];
                
                r_data[32936] <= r_data[32935];
                
                r_data[32937] <= r_data[32936];
                
                r_data[32938] <= r_data[32937];
                
                r_data[32939] <= r_data[32938];
                
                r_data[32940] <= r_data[32939];
                
                r_data[32941] <= r_data[32940];
                
                r_data[32942] <= r_data[32941];
                
                r_data[32943] <= r_data[32942];
                
                r_data[32944] <= r_data[32943];
                
                r_data[32945] <= r_data[32944];
                
                r_data[32946] <= r_data[32945];
                
                r_data[32947] <= r_data[32946];
                
                r_data[32948] <= r_data[32947];
                
                r_data[32949] <= r_data[32948];
                
                r_data[32950] <= r_data[32949];
                
                r_data[32951] <= r_data[32950];
                
                r_data[32952] <= r_data[32951];
                
                r_data[32953] <= r_data[32952];
                
                r_data[32954] <= r_data[32953];
                
                r_data[32955] <= r_data[32954];
                
                r_data[32956] <= r_data[32955];
                
                r_data[32957] <= r_data[32956];
                
                r_data[32958] <= r_data[32957];
                
                r_data[32959] <= r_data[32958];
                
                r_data[32960] <= r_data[32959];
                
                r_data[32961] <= r_data[32960];
                
                r_data[32962] <= r_data[32961];
                
                r_data[32963] <= r_data[32962];
                
                r_data[32964] <= r_data[32963];
                
                r_data[32965] <= r_data[32964];
                
                r_data[32966] <= r_data[32965];
                
                r_data[32967] <= r_data[32966];
                
                r_data[32968] <= r_data[32967];
                
                r_data[32969] <= r_data[32968];
                
                r_data[32970] <= r_data[32969];
                
                r_data[32971] <= r_data[32970];
                
                r_data[32972] <= r_data[32971];
                
                r_data[32973] <= r_data[32972];
                
                r_data[32974] <= r_data[32973];
                
                r_data[32975] <= r_data[32974];
                
                r_data[32976] <= r_data[32975];
                
                r_data[32977] <= r_data[32976];
                
                r_data[32978] <= r_data[32977];
                
                r_data[32979] <= r_data[32978];
                
                r_data[32980] <= r_data[32979];
                
                r_data[32981] <= r_data[32980];
                
                r_data[32982] <= r_data[32981];
                
                r_data[32983] <= r_data[32982];
                
                r_data[32984] <= r_data[32983];
                
                r_data[32985] <= r_data[32984];
                
                r_data[32986] <= r_data[32985];
                
                r_data[32987] <= r_data[32986];
                
                r_data[32988] <= r_data[32987];
                
                r_data[32989] <= r_data[32988];
                
                r_data[32990] <= r_data[32989];
                
                r_data[32991] <= r_data[32990];
                
                r_data[32992] <= r_data[32991];
                
                r_data[32993] <= r_data[32992];
                
                r_data[32994] <= r_data[32993];
                
                r_data[32995] <= r_data[32994];
                
                r_data[32996] <= r_data[32995];
                
                r_data[32997] <= r_data[32996];
                
                r_data[32998] <= r_data[32997];
                
                r_data[32999] <= r_data[32998];
                
                r_data[33000] <= r_data[32999];
                
                r_data[33001] <= r_data[33000];
                
                r_data[33002] <= r_data[33001];
                
                r_data[33003] <= r_data[33002];
                
                r_data[33004] <= r_data[33003];
                
                r_data[33005] <= r_data[33004];
                
                r_data[33006] <= r_data[33005];
                
                r_data[33007] <= r_data[33006];
                
                r_data[33008] <= r_data[33007];
                
                r_data[33009] <= r_data[33008];
                
                r_data[33010] <= r_data[33009];
                
                r_data[33011] <= r_data[33010];
                
                r_data[33012] <= r_data[33011];
                
                r_data[33013] <= r_data[33012];
                
                r_data[33014] <= r_data[33013];
                
                r_data[33015] <= r_data[33014];
                
                r_data[33016] <= r_data[33015];
                
                r_data[33017] <= r_data[33016];
                
                r_data[33018] <= r_data[33017];
                
                r_data[33019] <= r_data[33018];
                
                r_data[33020] <= r_data[33019];
                
                r_data[33021] <= r_data[33020];
                
                r_data[33022] <= r_data[33021];
                
                r_data[33023] <= r_data[33022];
                
                r_data[33024] <= r_data[33023];
                
                r_data[33025] <= r_data[33024];
                
                r_data[33026] <= r_data[33025];
                
                r_data[33027] <= r_data[33026];
                
                r_data[33028] <= r_data[33027];
                
                r_data[33029] <= r_data[33028];
                
                r_data[33030] <= r_data[33029];
                
                r_data[33031] <= r_data[33030];
                
                r_data[33032] <= r_data[33031];
                
                r_data[33033] <= r_data[33032];
                
                r_data[33034] <= r_data[33033];
                
                r_data[33035] <= r_data[33034];
                
                r_data[33036] <= r_data[33035];
                
                r_data[33037] <= r_data[33036];
                
                r_data[33038] <= r_data[33037];
                
                r_data[33039] <= r_data[33038];
                
                r_data[33040] <= r_data[33039];
                
                r_data[33041] <= r_data[33040];
                
                r_data[33042] <= r_data[33041];
                
                r_data[33043] <= r_data[33042];
                
                r_data[33044] <= r_data[33043];
                
                r_data[33045] <= r_data[33044];
                
                r_data[33046] <= r_data[33045];
                
                r_data[33047] <= r_data[33046];
                
                r_data[33048] <= r_data[33047];
                
                r_data[33049] <= r_data[33048];
                
                r_data[33050] <= r_data[33049];
                
                r_data[33051] <= r_data[33050];
                
                r_data[33052] <= r_data[33051];
                
                r_data[33053] <= r_data[33052];
                
                r_data[33054] <= r_data[33053];
                
                r_data[33055] <= r_data[33054];
                
                r_data[33056] <= r_data[33055];
                
                r_data[33057] <= r_data[33056];
                
                r_data[33058] <= r_data[33057];
                
                r_data[33059] <= r_data[33058];
                
                r_data[33060] <= r_data[33059];
                
                r_data[33061] <= r_data[33060];
                
                r_data[33062] <= r_data[33061];
                
                r_data[33063] <= r_data[33062];
                
                r_data[33064] <= r_data[33063];
                
                r_data[33065] <= r_data[33064];
                
                r_data[33066] <= r_data[33065];
                
                r_data[33067] <= r_data[33066];
                
                r_data[33068] <= r_data[33067];
                
                r_data[33069] <= r_data[33068];
                
                r_data[33070] <= r_data[33069];
                
                r_data[33071] <= r_data[33070];
                
                r_data[33072] <= r_data[33071];
                
                r_data[33073] <= r_data[33072];
                
                r_data[33074] <= r_data[33073];
                
                r_data[33075] <= r_data[33074];
                
                r_data[33076] <= r_data[33075];
                
                r_data[33077] <= r_data[33076];
                
                r_data[33078] <= r_data[33077];
                
                r_data[33079] <= r_data[33078];
                
                r_data[33080] <= r_data[33079];
                
                r_data[33081] <= r_data[33080];
                
                r_data[33082] <= r_data[33081];
                
                r_data[33083] <= r_data[33082];
                
                r_data[33084] <= r_data[33083];
                
                r_data[33085] <= r_data[33084];
                
                r_data[33086] <= r_data[33085];
                
                r_data[33087] <= r_data[33086];
                
                r_data[33088] <= r_data[33087];
                
                r_data[33089] <= r_data[33088];
                
                r_data[33090] <= r_data[33089];
                
                r_data[33091] <= r_data[33090];
                
                r_data[33092] <= r_data[33091];
                
                r_data[33093] <= r_data[33092];
                
                r_data[33094] <= r_data[33093];
                
                r_data[33095] <= r_data[33094];
                
                r_data[33096] <= r_data[33095];
                
                r_data[33097] <= r_data[33096];
                
                r_data[33098] <= r_data[33097];
                
                r_data[33099] <= r_data[33098];
                
                r_data[33100] <= r_data[33099];
                
                r_data[33101] <= r_data[33100];
                
                r_data[33102] <= r_data[33101];
                
                r_data[33103] <= r_data[33102];
                
                r_data[33104] <= r_data[33103];
                
                r_data[33105] <= r_data[33104];
                
                r_data[33106] <= r_data[33105];
                
                r_data[33107] <= r_data[33106];
                
                r_data[33108] <= r_data[33107];
                
                r_data[33109] <= r_data[33108];
                
                r_data[33110] <= r_data[33109];
                
                r_data[33111] <= r_data[33110];
                
                r_data[33112] <= r_data[33111];
                
                r_data[33113] <= r_data[33112];
                
                r_data[33114] <= r_data[33113];
                
                r_data[33115] <= r_data[33114];
                
                r_data[33116] <= r_data[33115];
                
                r_data[33117] <= r_data[33116];
                
                r_data[33118] <= r_data[33117];
                
                r_data[33119] <= r_data[33118];
                
                r_data[33120] <= r_data[33119];
                
                r_data[33121] <= r_data[33120];
                
                r_data[33122] <= r_data[33121];
                
                r_data[33123] <= r_data[33122];
                
                r_data[33124] <= r_data[33123];
                
                r_data[33125] <= r_data[33124];
                
                r_data[33126] <= r_data[33125];
                
                r_data[33127] <= r_data[33126];
                
                r_data[33128] <= r_data[33127];
                
                r_data[33129] <= r_data[33128];
                
                r_data[33130] <= r_data[33129];
                
                r_data[33131] <= r_data[33130];
                
                r_data[33132] <= r_data[33131];
                
                r_data[33133] <= r_data[33132];
                
                r_data[33134] <= r_data[33133];
                
                r_data[33135] <= r_data[33134];
                
                r_data[33136] <= r_data[33135];
                
                r_data[33137] <= r_data[33136];
                
                r_data[33138] <= r_data[33137];
                
                r_data[33139] <= r_data[33138];
                
                r_data[33140] <= r_data[33139];
                
                r_data[33141] <= r_data[33140];
                
                r_data[33142] <= r_data[33141];
                
                r_data[33143] <= r_data[33142];
                
                r_data[33144] <= r_data[33143];
                
                r_data[33145] <= r_data[33144];
                
                r_data[33146] <= r_data[33145];
                
                r_data[33147] <= r_data[33146];
                
                r_data[33148] <= r_data[33147];
                
                r_data[33149] <= r_data[33148];
                
                r_data[33150] <= r_data[33149];
                
                r_data[33151] <= r_data[33150];
                
                r_data[33152] <= r_data[33151];
                
                r_data[33153] <= r_data[33152];
                
                r_data[33154] <= r_data[33153];
                
                r_data[33155] <= r_data[33154];
                
                r_data[33156] <= r_data[33155];
                
                r_data[33157] <= r_data[33156];
                
                r_data[33158] <= r_data[33157];
                
                r_data[33159] <= r_data[33158];
                
                r_data[33160] <= r_data[33159];
                
                r_data[33161] <= r_data[33160];
                
                r_data[33162] <= r_data[33161];
                
                r_data[33163] <= r_data[33162];
                
                r_data[33164] <= r_data[33163];
                
                r_data[33165] <= r_data[33164];
                
                r_data[33166] <= r_data[33165];
                
                r_data[33167] <= r_data[33166];
                
                r_data[33168] <= r_data[33167];
                
                r_data[33169] <= r_data[33168];
                
                r_data[33170] <= r_data[33169];
                
                r_data[33171] <= r_data[33170];
                
                r_data[33172] <= r_data[33171];
                
                r_data[33173] <= r_data[33172];
                
                r_data[33174] <= r_data[33173];
                
                r_data[33175] <= r_data[33174];
                
                r_data[33176] <= r_data[33175];
                
                r_data[33177] <= r_data[33176];
                
                r_data[33178] <= r_data[33177];
                
                r_data[33179] <= r_data[33178];
                
                r_data[33180] <= r_data[33179];
                
                r_data[33181] <= r_data[33180];
                
                r_data[33182] <= r_data[33181];
                
                r_data[33183] <= r_data[33182];
                
                r_data[33184] <= r_data[33183];
                
                r_data[33185] <= r_data[33184];
                
                r_data[33186] <= r_data[33185];
                
                r_data[33187] <= r_data[33186];
                
                r_data[33188] <= r_data[33187];
                
                r_data[33189] <= r_data[33188];
                
                r_data[33190] <= r_data[33189];
                
                r_data[33191] <= r_data[33190];
                
                r_data[33192] <= r_data[33191];
                
                r_data[33193] <= r_data[33192];
                
                r_data[33194] <= r_data[33193];
                
                r_data[33195] <= r_data[33194];
                
                r_data[33196] <= r_data[33195];
                
                r_data[33197] <= r_data[33196];
                
                r_data[33198] <= r_data[33197];
                
                r_data[33199] <= r_data[33198];
                
                r_data[33200] <= r_data[33199];
                
                r_data[33201] <= r_data[33200];
                
                r_data[33202] <= r_data[33201];
                
                r_data[33203] <= r_data[33202];
                
                r_data[33204] <= r_data[33203];
                
                r_data[33205] <= r_data[33204];
                
                r_data[33206] <= r_data[33205];
                
                r_data[33207] <= r_data[33206];
                
                r_data[33208] <= r_data[33207];
                
                r_data[33209] <= r_data[33208];
                
                r_data[33210] <= r_data[33209];
                
                r_data[33211] <= r_data[33210];
                
                r_data[33212] <= r_data[33211];
                
                r_data[33213] <= r_data[33212];
                
                r_data[33214] <= r_data[33213];
                
                r_data[33215] <= r_data[33214];
                
                r_data[33216] <= r_data[33215];
                
                r_data[33217] <= r_data[33216];
                
                r_data[33218] <= r_data[33217];
                
                r_data[33219] <= r_data[33218];
                
                r_data[33220] <= r_data[33219];
                
                r_data[33221] <= r_data[33220];
                
                r_data[33222] <= r_data[33221];
                
                r_data[33223] <= r_data[33222];
                
                r_data[33224] <= r_data[33223];
                
                r_data[33225] <= r_data[33224];
                
                r_data[33226] <= r_data[33225];
                
                r_data[33227] <= r_data[33226];
                
                r_data[33228] <= r_data[33227];
                
                r_data[33229] <= r_data[33228];
                
                r_data[33230] <= r_data[33229];
                
                r_data[33231] <= r_data[33230];
                
                r_data[33232] <= r_data[33231];
                
                r_data[33233] <= r_data[33232];
                
                r_data[33234] <= r_data[33233];
                
                r_data[33235] <= r_data[33234];
                
                r_data[33236] <= r_data[33235];
                
                r_data[33237] <= r_data[33236];
                
                r_data[33238] <= r_data[33237];
                
                r_data[33239] <= r_data[33238];
                
                r_data[33240] <= r_data[33239];
                
                r_data[33241] <= r_data[33240];
                
                r_data[33242] <= r_data[33241];
                
                r_data[33243] <= r_data[33242];
                
                r_data[33244] <= r_data[33243];
                
                r_data[33245] <= r_data[33244];
                
                r_data[33246] <= r_data[33245];
                
                r_data[33247] <= r_data[33246];
                
                r_data[33248] <= r_data[33247];
                
                r_data[33249] <= r_data[33248];
                
                r_data[33250] <= r_data[33249];
                
                r_data[33251] <= r_data[33250];
                
                r_data[33252] <= r_data[33251];
                
                r_data[33253] <= r_data[33252];
                
                r_data[33254] <= r_data[33253];
                
                r_data[33255] <= r_data[33254];
                
                r_data[33256] <= r_data[33255];
                
                r_data[33257] <= r_data[33256];
                
                r_data[33258] <= r_data[33257];
                
                r_data[33259] <= r_data[33258];
                
                r_data[33260] <= r_data[33259];
                
                r_data[33261] <= r_data[33260];
                
                r_data[33262] <= r_data[33261];
                
                r_data[33263] <= r_data[33262];
                
                r_data[33264] <= r_data[33263];
                
                r_data[33265] <= r_data[33264];
                
                r_data[33266] <= r_data[33265];
                
                r_data[33267] <= r_data[33266];
                
                r_data[33268] <= r_data[33267];
                
                r_data[33269] <= r_data[33268];
                
                r_data[33270] <= r_data[33269];
                
                r_data[33271] <= r_data[33270];
                
                r_data[33272] <= r_data[33271];
                
                r_data[33273] <= r_data[33272];
                
                r_data[33274] <= r_data[33273];
                
                r_data[33275] <= r_data[33274];
                
                r_data[33276] <= r_data[33275];
                
                r_data[33277] <= r_data[33276];
                
                r_data[33278] <= r_data[33277];
                
                r_data[33279] <= r_data[33278];
                
                r_data[33280] <= r_data[33279];
                
                r_data[33281] <= r_data[33280];
                
                r_data[33282] <= r_data[33281];
                
                r_data[33283] <= r_data[33282];
                
                r_data[33284] <= r_data[33283];
                
                r_data[33285] <= r_data[33284];
                
                r_data[33286] <= r_data[33285];
                
                r_data[33287] <= r_data[33286];
                
                r_data[33288] <= r_data[33287];
                
                r_data[33289] <= r_data[33288];
                
                r_data[33290] <= r_data[33289];
                
                r_data[33291] <= r_data[33290];
                
                r_data[33292] <= r_data[33291];
                
                r_data[33293] <= r_data[33292];
                
                r_data[33294] <= r_data[33293];
                
                r_data[33295] <= r_data[33294];
                
                r_data[33296] <= r_data[33295];
                
                r_data[33297] <= r_data[33296];
                
                r_data[33298] <= r_data[33297];
                
                r_data[33299] <= r_data[33298];
                
                r_data[33300] <= r_data[33299];
                
                r_data[33301] <= r_data[33300];
                
                r_data[33302] <= r_data[33301];
                
                r_data[33303] <= r_data[33302];
                
                r_data[33304] <= r_data[33303];
                
                r_data[33305] <= r_data[33304];
                
                r_data[33306] <= r_data[33305];
                
                r_data[33307] <= r_data[33306];
                
                r_data[33308] <= r_data[33307];
                
                r_data[33309] <= r_data[33308];
                
                r_data[33310] <= r_data[33309];
                
                r_data[33311] <= r_data[33310];
                
                r_data[33312] <= r_data[33311];
                
                r_data[33313] <= r_data[33312];
                
                r_data[33314] <= r_data[33313];
                
                r_data[33315] <= r_data[33314];
                
                r_data[33316] <= r_data[33315];
                
                r_data[33317] <= r_data[33316];
                
                r_data[33318] <= r_data[33317];
                
                r_data[33319] <= r_data[33318];
                
                r_data[33320] <= r_data[33319];
                
                r_data[33321] <= r_data[33320];
                
                r_data[33322] <= r_data[33321];
                
                r_data[33323] <= r_data[33322];
                
                r_data[33324] <= r_data[33323];
                
                r_data[33325] <= r_data[33324];
                
                r_data[33326] <= r_data[33325];
                
                r_data[33327] <= r_data[33326];
                
                r_data[33328] <= r_data[33327];
                
                r_data[33329] <= r_data[33328];
                
                r_data[33330] <= r_data[33329];
                
                r_data[33331] <= r_data[33330];
                
                r_data[33332] <= r_data[33331];
                
                r_data[33333] <= r_data[33332];
                
                r_data[33334] <= r_data[33333];
                
                r_data[33335] <= r_data[33334];
                
                r_data[33336] <= r_data[33335];
                
                r_data[33337] <= r_data[33336];
                
                r_data[33338] <= r_data[33337];
                
                r_data[33339] <= r_data[33338];
                
                r_data[33340] <= r_data[33339];
                
                r_data[33341] <= r_data[33340];
                
                r_data[33342] <= r_data[33341];
                
                r_data[33343] <= r_data[33342];
                
                r_data[33344] <= r_data[33343];
                
                r_data[33345] <= r_data[33344];
                
                r_data[33346] <= r_data[33345];
                
                r_data[33347] <= r_data[33346];
                
                r_data[33348] <= r_data[33347];
                
                r_data[33349] <= r_data[33348];
                
                r_data[33350] <= r_data[33349];
                
                r_data[33351] <= r_data[33350];
                
                r_data[33352] <= r_data[33351];
                
                r_data[33353] <= r_data[33352];
                
                r_data[33354] <= r_data[33353];
                
                r_data[33355] <= r_data[33354];
                
                r_data[33356] <= r_data[33355];
                
                r_data[33357] <= r_data[33356];
                
                r_data[33358] <= r_data[33357];
                
                r_data[33359] <= r_data[33358];
                
                r_data[33360] <= r_data[33359];
                
                r_data[33361] <= r_data[33360];
                
                r_data[33362] <= r_data[33361];
                
                r_data[33363] <= r_data[33362];
                
                r_data[33364] <= r_data[33363];
                
                r_data[33365] <= r_data[33364];
                
                r_data[33366] <= r_data[33365];
                
                r_data[33367] <= r_data[33366];
                
                r_data[33368] <= r_data[33367];
                
                r_data[33369] <= r_data[33368];
                
                r_data[33370] <= r_data[33369];
                
                r_data[33371] <= r_data[33370];
                
                r_data[33372] <= r_data[33371];
                
                r_data[33373] <= r_data[33372];
                
                r_data[33374] <= r_data[33373];
                
                r_data[33375] <= r_data[33374];
                
                r_data[33376] <= r_data[33375];
                
                r_data[33377] <= r_data[33376];
                
                r_data[33378] <= r_data[33377];
                
                r_data[33379] <= r_data[33378];
                
                r_data[33380] <= r_data[33379];
                
                r_data[33381] <= r_data[33380];
                
                r_data[33382] <= r_data[33381];
                
                r_data[33383] <= r_data[33382];
                
                r_data[33384] <= r_data[33383];
                
                r_data[33385] <= r_data[33384];
                
                r_data[33386] <= r_data[33385];
                
                r_data[33387] <= r_data[33386];
                
                r_data[33388] <= r_data[33387];
                
                r_data[33389] <= r_data[33388];
                
                r_data[33390] <= r_data[33389];
                
                r_data[33391] <= r_data[33390];
                
                r_data[33392] <= r_data[33391];
                
                r_data[33393] <= r_data[33392];
                
                r_data[33394] <= r_data[33393];
                
                r_data[33395] <= r_data[33394];
                
                r_data[33396] <= r_data[33395];
                
                r_data[33397] <= r_data[33396];
                
                r_data[33398] <= r_data[33397];
                
                r_data[33399] <= r_data[33398];
                
                r_data[33400] <= r_data[33399];
                
                r_data[33401] <= r_data[33400];
                
                r_data[33402] <= r_data[33401];
                
                r_data[33403] <= r_data[33402];
                
                r_data[33404] <= r_data[33403];
                
                r_data[33405] <= r_data[33404];
                
                r_data[33406] <= r_data[33405];
                
                r_data[33407] <= r_data[33406];
                
                r_data[33408] <= r_data[33407];
                
                r_data[33409] <= r_data[33408];
                
                r_data[33410] <= r_data[33409];
                
                r_data[33411] <= r_data[33410];
                
                r_data[33412] <= r_data[33411];
                
                r_data[33413] <= r_data[33412];
                
                r_data[33414] <= r_data[33413];
                
                r_data[33415] <= r_data[33414];
                
                r_data[33416] <= r_data[33415];
                
                r_data[33417] <= r_data[33416];
                
                r_data[33418] <= r_data[33417];
                
                r_data[33419] <= r_data[33418];
                
                r_data[33420] <= r_data[33419];
                
                r_data[33421] <= r_data[33420];
                
                r_data[33422] <= r_data[33421];
                
                r_data[33423] <= r_data[33422];
                
                r_data[33424] <= r_data[33423];
                
                r_data[33425] <= r_data[33424];
                
                r_data[33426] <= r_data[33425];
                
                r_data[33427] <= r_data[33426];
                
                r_data[33428] <= r_data[33427];
                
                r_data[33429] <= r_data[33428];
                
                r_data[33430] <= r_data[33429];
                
                r_data[33431] <= r_data[33430];
                
                r_data[33432] <= r_data[33431];
                
                r_data[33433] <= r_data[33432];
                
                r_data[33434] <= r_data[33433];
                
                r_data[33435] <= r_data[33434];
                
                r_data[33436] <= r_data[33435];
                
                r_data[33437] <= r_data[33436];
                
                r_data[33438] <= r_data[33437];
                
                r_data[33439] <= r_data[33438];
                
                r_data[33440] <= r_data[33439];
                
                r_data[33441] <= r_data[33440];
                
                r_data[33442] <= r_data[33441];
                
                r_data[33443] <= r_data[33442];
                
                r_data[33444] <= r_data[33443];
                
                r_data[33445] <= r_data[33444];
                
                r_data[33446] <= r_data[33445];
                
                r_data[33447] <= r_data[33446];
                
                r_data[33448] <= r_data[33447];
                
                r_data[33449] <= r_data[33448];
                
                r_data[33450] <= r_data[33449];
                
                r_data[33451] <= r_data[33450];
                
                r_data[33452] <= r_data[33451];
                
                r_data[33453] <= r_data[33452];
                
                r_data[33454] <= r_data[33453];
                
                r_data[33455] <= r_data[33454];
                
                r_data[33456] <= r_data[33455];
                
                r_data[33457] <= r_data[33456];
                
                r_data[33458] <= r_data[33457];
                
                r_data[33459] <= r_data[33458];
                
                r_data[33460] <= r_data[33459];
                
                r_data[33461] <= r_data[33460];
                
                r_data[33462] <= r_data[33461];
                
                r_data[33463] <= r_data[33462];
                
                r_data[33464] <= r_data[33463];
                
                r_data[33465] <= r_data[33464];
                
                r_data[33466] <= r_data[33465];
                
                r_data[33467] <= r_data[33466];
                
                r_data[33468] <= r_data[33467];
                
                r_data[33469] <= r_data[33468];
                
                r_data[33470] <= r_data[33469];
                
                r_data[33471] <= r_data[33470];
                
                r_data[33472] <= r_data[33471];
                
                r_data[33473] <= r_data[33472];
                
                r_data[33474] <= r_data[33473];
                
                r_data[33475] <= r_data[33474];
                
                r_data[33476] <= r_data[33475];
                
                r_data[33477] <= r_data[33476];
                
                r_data[33478] <= r_data[33477];
                
                r_data[33479] <= r_data[33478];
                
                r_data[33480] <= r_data[33479];
                
                r_data[33481] <= r_data[33480];
                
                r_data[33482] <= r_data[33481];
                
                r_data[33483] <= r_data[33482];
                
                r_data[33484] <= r_data[33483];
                
                r_data[33485] <= r_data[33484];
                
                r_data[33486] <= r_data[33485];
                
                r_data[33487] <= r_data[33486];
                
                r_data[33488] <= r_data[33487];
                
                r_data[33489] <= r_data[33488];
                
                r_data[33490] <= r_data[33489];
                
                r_data[33491] <= r_data[33490];
                
                r_data[33492] <= r_data[33491];
                
                r_data[33493] <= r_data[33492];
                
                r_data[33494] <= r_data[33493];
                
                r_data[33495] <= r_data[33494];
                
                r_data[33496] <= r_data[33495];
                
                r_data[33497] <= r_data[33496];
                
                r_data[33498] <= r_data[33497];
                
                r_data[33499] <= r_data[33498];
                
                r_data[33500] <= r_data[33499];
                
                r_data[33501] <= r_data[33500];
                
                r_data[33502] <= r_data[33501];
                
                r_data[33503] <= r_data[33502];
                
                r_data[33504] <= r_data[33503];
                
                r_data[33505] <= r_data[33504];
                
                r_data[33506] <= r_data[33505];
                
                r_data[33507] <= r_data[33506];
                
                r_data[33508] <= r_data[33507];
                
                r_data[33509] <= r_data[33508];
                
                r_data[33510] <= r_data[33509];
                
                r_data[33511] <= r_data[33510];
                
                r_data[33512] <= r_data[33511];
                
                r_data[33513] <= r_data[33512];
                
                r_data[33514] <= r_data[33513];
                
                r_data[33515] <= r_data[33514];
                
                r_data[33516] <= r_data[33515];
                
                r_data[33517] <= r_data[33516];
                
                r_data[33518] <= r_data[33517];
                
                r_data[33519] <= r_data[33518];
                
                r_data[33520] <= r_data[33519];
                
                r_data[33521] <= r_data[33520];
                
                r_data[33522] <= r_data[33521];
                
                r_data[33523] <= r_data[33522];
                
                r_data[33524] <= r_data[33523];
                
                r_data[33525] <= r_data[33524];
                
                r_data[33526] <= r_data[33525];
                
                r_data[33527] <= r_data[33526];
                
                r_data[33528] <= r_data[33527];
                
                r_data[33529] <= r_data[33528];
                
                r_data[33530] <= r_data[33529];
                
                r_data[33531] <= r_data[33530];
                
                r_data[33532] <= r_data[33531];
                
                r_data[33533] <= r_data[33532];
                
                r_data[33534] <= r_data[33533];
                
                r_data[33535] <= r_data[33534];
                
                r_data[33536] <= r_data[33535];
                
                r_data[33537] <= r_data[33536];
                
                r_data[33538] <= r_data[33537];
                
                r_data[33539] <= r_data[33538];
                
                r_data[33540] <= r_data[33539];
                
                r_data[33541] <= r_data[33540];
                
                r_data[33542] <= r_data[33541];
                
                r_data[33543] <= r_data[33542];
                
                r_data[33544] <= r_data[33543];
                
                r_data[33545] <= r_data[33544];
                
                r_data[33546] <= r_data[33545];
                
                r_data[33547] <= r_data[33546];
                
                r_data[33548] <= r_data[33547];
                
                r_data[33549] <= r_data[33548];
                
                r_data[33550] <= r_data[33549];
                
                r_data[33551] <= r_data[33550];
                
                r_data[33552] <= r_data[33551];
                
                r_data[33553] <= r_data[33552];
                
                r_data[33554] <= r_data[33553];
                
                r_data[33555] <= r_data[33554];
                
                r_data[33556] <= r_data[33555];
                
                r_data[33557] <= r_data[33556];
                
                r_data[33558] <= r_data[33557];
                
                r_data[33559] <= r_data[33558];
                
                r_data[33560] <= r_data[33559];
                
                r_data[33561] <= r_data[33560];
                
                r_data[33562] <= r_data[33561];
                
                r_data[33563] <= r_data[33562];
                
                r_data[33564] <= r_data[33563];
                
                r_data[33565] <= r_data[33564];
                
                r_data[33566] <= r_data[33565];
                
                r_data[33567] <= r_data[33566];
                
                r_data[33568] <= r_data[33567];
                
                r_data[33569] <= r_data[33568];
                
                r_data[33570] <= r_data[33569];
                
                r_data[33571] <= r_data[33570];
                
                r_data[33572] <= r_data[33571];
                
                r_data[33573] <= r_data[33572];
                
                r_data[33574] <= r_data[33573];
                
                r_data[33575] <= r_data[33574];
                
                r_data[33576] <= r_data[33575];
                
                r_data[33577] <= r_data[33576];
                
                r_data[33578] <= r_data[33577];
                
                r_data[33579] <= r_data[33578];
                
                r_data[33580] <= r_data[33579];
                
                r_data[33581] <= r_data[33580];
                
                r_data[33582] <= r_data[33581];
                
                r_data[33583] <= r_data[33582];
                
                r_data[33584] <= r_data[33583];
                
                r_data[33585] <= r_data[33584];
                
                r_data[33586] <= r_data[33585];
                
                r_data[33587] <= r_data[33586];
                
                r_data[33588] <= r_data[33587];
                
                r_data[33589] <= r_data[33588];
                
                r_data[33590] <= r_data[33589];
                
                r_data[33591] <= r_data[33590];
                
                r_data[33592] <= r_data[33591];
                
                r_data[33593] <= r_data[33592];
                
                r_data[33594] <= r_data[33593];
                
                r_data[33595] <= r_data[33594];
                
                r_data[33596] <= r_data[33595];
                
                r_data[33597] <= r_data[33596];
                
                r_data[33598] <= r_data[33597];
                
                r_data[33599] <= r_data[33598];
                
                r_data[33600] <= r_data[33599];
                
                r_data[33601] <= r_data[33600];
                
                r_data[33602] <= r_data[33601];
                
                r_data[33603] <= r_data[33602];
                
                r_data[33604] <= r_data[33603];
                
                r_data[33605] <= r_data[33604];
                
                r_data[33606] <= r_data[33605];
                
                r_data[33607] <= r_data[33606];
                
                r_data[33608] <= r_data[33607];
                
                r_data[33609] <= r_data[33608];
                
                r_data[33610] <= r_data[33609];
                
                r_data[33611] <= r_data[33610];
                
                r_data[33612] <= r_data[33611];
                
                r_data[33613] <= r_data[33612];
                
                r_data[33614] <= r_data[33613];
                
                r_data[33615] <= r_data[33614];
                
                r_data[33616] <= r_data[33615];
                
                r_data[33617] <= r_data[33616];
                
                r_data[33618] <= r_data[33617];
                
                r_data[33619] <= r_data[33618];
                
                r_data[33620] <= r_data[33619];
                
                r_data[33621] <= r_data[33620];
                
                r_data[33622] <= r_data[33621];
                
                r_data[33623] <= r_data[33622];
                
                r_data[33624] <= r_data[33623];
                
                r_data[33625] <= r_data[33624];
                
                r_data[33626] <= r_data[33625];
                
                r_data[33627] <= r_data[33626];
                
                r_data[33628] <= r_data[33627];
                
                r_data[33629] <= r_data[33628];
                
                r_data[33630] <= r_data[33629];
                
                r_data[33631] <= r_data[33630];
                
                r_data[33632] <= r_data[33631];
                
                r_data[33633] <= r_data[33632];
                
                r_data[33634] <= r_data[33633];
                
                r_data[33635] <= r_data[33634];
                
                r_data[33636] <= r_data[33635];
                
                r_data[33637] <= r_data[33636];
                
                r_data[33638] <= r_data[33637];
                
                r_data[33639] <= r_data[33638];
                
                r_data[33640] <= r_data[33639];
                
                r_data[33641] <= r_data[33640];
                
                r_data[33642] <= r_data[33641];
                
                r_data[33643] <= r_data[33642];
                
                r_data[33644] <= r_data[33643];
                
                r_data[33645] <= r_data[33644];
                
                r_data[33646] <= r_data[33645];
                
                r_data[33647] <= r_data[33646];
                
                r_data[33648] <= r_data[33647];
                
                r_data[33649] <= r_data[33648];
                
                r_data[33650] <= r_data[33649];
                
                r_data[33651] <= r_data[33650];
                
                r_data[33652] <= r_data[33651];
                
                r_data[33653] <= r_data[33652];
                
                r_data[33654] <= r_data[33653];
                
                r_data[33655] <= r_data[33654];
                
                r_data[33656] <= r_data[33655];
                
                r_data[33657] <= r_data[33656];
                
                r_data[33658] <= r_data[33657];
                
                r_data[33659] <= r_data[33658];
                
                r_data[33660] <= r_data[33659];
                
                r_data[33661] <= r_data[33660];
                
                r_data[33662] <= r_data[33661];
                
                r_data[33663] <= r_data[33662];
                
                r_data[33664] <= r_data[33663];
                
                r_data[33665] <= r_data[33664];
                
                r_data[33666] <= r_data[33665];
                
                r_data[33667] <= r_data[33666];
                
                r_data[33668] <= r_data[33667];
                
                r_data[33669] <= r_data[33668];
                
                r_data[33670] <= r_data[33669];
                
                r_data[33671] <= r_data[33670];
                
                r_data[33672] <= r_data[33671];
                
                r_data[33673] <= r_data[33672];
                
                r_data[33674] <= r_data[33673];
                
                r_data[33675] <= r_data[33674];
                
                r_data[33676] <= r_data[33675];
                
                r_data[33677] <= r_data[33676];
                
                r_data[33678] <= r_data[33677];
                
                r_data[33679] <= r_data[33678];
                
                r_data[33680] <= r_data[33679];
                
                r_data[33681] <= r_data[33680];
                
                r_data[33682] <= r_data[33681];
                
                r_data[33683] <= r_data[33682];
                
                r_data[33684] <= r_data[33683];
                
                r_data[33685] <= r_data[33684];
                
                r_data[33686] <= r_data[33685];
                
                r_data[33687] <= r_data[33686];
                
                r_data[33688] <= r_data[33687];
                
                r_data[33689] <= r_data[33688];
                
                r_data[33690] <= r_data[33689];
                
                r_data[33691] <= r_data[33690];
                
                r_data[33692] <= r_data[33691];
                
                r_data[33693] <= r_data[33692];
                
                r_data[33694] <= r_data[33693];
                
                r_data[33695] <= r_data[33694];
                
                r_data[33696] <= r_data[33695];
                
                r_data[33697] <= r_data[33696];
                
                r_data[33698] <= r_data[33697];
                
                r_data[33699] <= r_data[33698];
                
                r_data[33700] <= r_data[33699];
                
                r_data[33701] <= r_data[33700];
                
                r_data[33702] <= r_data[33701];
                
                r_data[33703] <= r_data[33702];
                
                r_data[33704] <= r_data[33703];
                
                r_data[33705] <= r_data[33704];
                
                r_data[33706] <= r_data[33705];
                
                r_data[33707] <= r_data[33706];
                
                r_data[33708] <= r_data[33707];
                
                r_data[33709] <= r_data[33708];
                
                r_data[33710] <= r_data[33709];
                
                r_data[33711] <= r_data[33710];
                
                r_data[33712] <= r_data[33711];
                
                r_data[33713] <= r_data[33712];
                
                r_data[33714] <= r_data[33713];
                
                r_data[33715] <= r_data[33714];
                
                r_data[33716] <= r_data[33715];
                
                r_data[33717] <= r_data[33716];
                
                r_data[33718] <= r_data[33717];
                
                r_data[33719] <= r_data[33718];
                
                r_data[33720] <= r_data[33719];
                
                r_data[33721] <= r_data[33720];
                
                r_data[33722] <= r_data[33721];
                
                r_data[33723] <= r_data[33722];
                
                r_data[33724] <= r_data[33723];
                
                r_data[33725] <= r_data[33724];
                
                r_data[33726] <= r_data[33725];
                
                r_data[33727] <= r_data[33726];
                
                r_data[33728] <= r_data[33727];
                
                r_data[33729] <= r_data[33728];
                
                r_data[33730] <= r_data[33729];
                
                r_data[33731] <= r_data[33730];
                
                r_data[33732] <= r_data[33731];
                
                r_data[33733] <= r_data[33732];
                
                r_data[33734] <= r_data[33733];
                
                r_data[33735] <= r_data[33734];
                
                r_data[33736] <= r_data[33735];
                
                r_data[33737] <= r_data[33736];
                
                r_data[33738] <= r_data[33737];
                
                r_data[33739] <= r_data[33738];
                
                r_data[33740] <= r_data[33739];
                
                r_data[33741] <= r_data[33740];
                
                r_data[33742] <= r_data[33741];
                
                r_data[33743] <= r_data[33742];
                
                r_data[33744] <= r_data[33743];
                
                r_data[33745] <= r_data[33744];
                
                r_data[33746] <= r_data[33745];
                
                r_data[33747] <= r_data[33746];
                
                r_data[33748] <= r_data[33747];
                
                r_data[33749] <= r_data[33748];
                
                r_data[33750] <= r_data[33749];
                
                r_data[33751] <= r_data[33750];
                
                r_data[33752] <= r_data[33751];
                
                r_data[33753] <= r_data[33752];
                
                r_data[33754] <= r_data[33753];
                
                r_data[33755] <= r_data[33754];
                
                r_data[33756] <= r_data[33755];
                
                r_data[33757] <= r_data[33756];
                
                r_data[33758] <= r_data[33757];
                
                r_data[33759] <= r_data[33758];
                
                r_data[33760] <= r_data[33759];
                
                r_data[33761] <= r_data[33760];
                
                r_data[33762] <= r_data[33761];
                
                r_data[33763] <= r_data[33762];
                
                r_data[33764] <= r_data[33763];
                
                r_data[33765] <= r_data[33764];
                
                r_data[33766] <= r_data[33765];
                
                r_data[33767] <= r_data[33766];
                
                r_data[33768] <= r_data[33767];
                
                r_data[33769] <= r_data[33768];
                
                r_data[33770] <= r_data[33769];
                
                r_data[33771] <= r_data[33770];
                
                r_data[33772] <= r_data[33771];
                
                r_data[33773] <= r_data[33772];
                
                r_data[33774] <= r_data[33773];
                
                r_data[33775] <= r_data[33774];
                
                r_data[33776] <= r_data[33775];
                
                r_data[33777] <= r_data[33776];
                
                r_data[33778] <= r_data[33777];
                
                r_data[33779] <= r_data[33778];
                
                r_data[33780] <= r_data[33779];
                
                r_data[33781] <= r_data[33780];
                
                r_data[33782] <= r_data[33781];
                
                r_data[33783] <= r_data[33782];
                
                r_data[33784] <= r_data[33783];
                
                r_data[33785] <= r_data[33784];
                
                r_data[33786] <= r_data[33785];
                
                r_data[33787] <= r_data[33786];
                
                r_data[33788] <= r_data[33787];
                
                r_data[33789] <= r_data[33788];
                
                r_data[33790] <= r_data[33789];
                
                r_data[33791] <= r_data[33790];
                
                r_data[33792] <= r_data[33791];
                
                r_data[33793] <= r_data[33792];
                
                r_data[33794] <= r_data[33793];
                
                r_data[33795] <= r_data[33794];
                
                r_data[33796] <= r_data[33795];
                
                r_data[33797] <= r_data[33796];
                
                r_data[33798] <= r_data[33797];
                
                r_data[33799] <= r_data[33798];
                
                r_data[33800] <= r_data[33799];
                
                r_data[33801] <= r_data[33800];
                
                r_data[33802] <= r_data[33801];
                
                r_data[33803] <= r_data[33802];
                
                r_data[33804] <= r_data[33803];
                
                r_data[33805] <= r_data[33804];
                
                r_data[33806] <= r_data[33805];
                
                r_data[33807] <= r_data[33806];
                
                r_data[33808] <= r_data[33807];
                
                r_data[33809] <= r_data[33808];
                
                r_data[33810] <= r_data[33809];
                
                r_data[33811] <= r_data[33810];
                
                r_data[33812] <= r_data[33811];
                
                r_data[33813] <= r_data[33812];
                
                r_data[33814] <= r_data[33813];
                
                r_data[33815] <= r_data[33814];
                
                r_data[33816] <= r_data[33815];
                
                r_data[33817] <= r_data[33816];
                
                r_data[33818] <= r_data[33817];
                
                r_data[33819] <= r_data[33818];
                
                r_data[33820] <= r_data[33819];
                
                r_data[33821] <= r_data[33820];
                
                r_data[33822] <= r_data[33821];
                
                r_data[33823] <= r_data[33822];
                
                r_data[33824] <= r_data[33823];
                
                r_data[33825] <= r_data[33824];
                
                r_data[33826] <= r_data[33825];
                
                r_data[33827] <= r_data[33826];
                
                r_data[33828] <= r_data[33827];
                
                r_data[33829] <= r_data[33828];
                
                r_data[33830] <= r_data[33829];
                
                r_data[33831] <= r_data[33830];
                
                r_data[33832] <= r_data[33831];
                
                r_data[33833] <= r_data[33832];
                
                r_data[33834] <= r_data[33833];
                
                r_data[33835] <= r_data[33834];
                
                r_data[33836] <= r_data[33835];
                
                r_data[33837] <= r_data[33836];
                
                r_data[33838] <= r_data[33837];
                
                r_data[33839] <= r_data[33838];
                
                r_data[33840] <= r_data[33839];
                
                r_data[33841] <= r_data[33840];
                
                r_data[33842] <= r_data[33841];
                
                r_data[33843] <= r_data[33842];
                
                r_data[33844] <= r_data[33843];
                
                r_data[33845] <= r_data[33844];
                
                r_data[33846] <= r_data[33845];
                
                r_data[33847] <= r_data[33846];
                
                r_data[33848] <= r_data[33847];
                
                r_data[33849] <= r_data[33848];
                
                r_data[33850] <= r_data[33849];
                
                r_data[33851] <= r_data[33850];
                
                r_data[33852] <= r_data[33851];
                
                r_data[33853] <= r_data[33852];
                
                r_data[33854] <= r_data[33853];
                
                r_data[33855] <= r_data[33854];
                
                r_data[33856] <= r_data[33855];
                
                r_data[33857] <= r_data[33856];
                
                r_data[33858] <= r_data[33857];
                
                r_data[33859] <= r_data[33858];
                
                r_data[33860] <= r_data[33859];
                
                r_data[33861] <= r_data[33860];
                
                r_data[33862] <= r_data[33861];
                
                r_data[33863] <= r_data[33862];
                
                r_data[33864] <= r_data[33863];
                
                r_data[33865] <= r_data[33864];
                
                r_data[33866] <= r_data[33865];
                
                r_data[33867] <= r_data[33866];
                
                r_data[33868] <= r_data[33867];
                
                r_data[33869] <= r_data[33868];
                
                r_data[33870] <= r_data[33869];
                
                r_data[33871] <= r_data[33870];
                
                r_data[33872] <= r_data[33871];
                
                r_data[33873] <= r_data[33872];
                
                r_data[33874] <= r_data[33873];
                
                r_data[33875] <= r_data[33874];
                
                r_data[33876] <= r_data[33875];
                
                r_data[33877] <= r_data[33876];
                
                r_data[33878] <= r_data[33877];
                
                r_data[33879] <= r_data[33878];
                
                r_data[33880] <= r_data[33879];
                
                r_data[33881] <= r_data[33880];
                
                r_data[33882] <= r_data[33881];
                
                r_data[33883] <= r_data[33882];
                
                r_data[33884] <= r_data[33883];
                
                r_data[33885] <= r_data[33884];
                
                r_data[33886] <= r_data[33885];
                
                r_data[33887] <= r_data[33886];
                
                r_data[33888] <= r_data[33887];
                
                r_data[33889] <= r_data[33888];
                
                r_data[33890] <= r_data[33889];
                
                r_data[33891] <= r_data[33890];
                
                r_data[33892] <= r_data[33891];
                
                r_data[33893] <= r_data[33892];
                
                r_data[33894] <= r_data[33893];
                
                r_data[33895] <= r_data[33894];
                
                r_data[33896] <= r_data[33895];
                
                r_data[33897] <= r_data[33896];
                
                r_data[33898] <= r_data[33897];
                
                r_data[33899] <= r_data[33898];
                
                r_data[33900] <= r_data[33899];
                
                r_data[33901] <= r_data[33900];
                
                r_data[33902] <= r_data[33901];
                
                r_data[33903] <= r_data[33902];
                
                r_data[33904] <= r_data[33903];
                
                r_data[33905] <= r_data[33904];
                
                r_data[33906] <= r_data[33905];
                
                r_data[33907] <= r_data[33906];
                
                r_data[33908] <= r_data[33907];
                
                r_data[33909] <= r_data[33908];
                
                r_data[33910] <= r_data[33909];
                
                r_data[33911] <= r_data[33910];
                
                r_data[33912] <= r_data[33911];
                
                r_data[33913] <= r_data[33912];
                
                r_data[33914] <= r_data[33913];
                
                r_data[33915] <= r_data[33914];
                
                r_data[33916] <= r_data[33915];
                
                r_data[33917] <= r_data[33916];
                
                r_data[33918] <= r_data[33917];
                
                r_data[33919] <= r_data[33918];
                
                r_data[33920] <= r_data[33919];
                
                r_data[33921] <= r_data[33920];
                
                r_data[33922] <= r_data[33921];
                
                r_data[33923] <= r_data[33922];
                
                r_data[33924] <= r_data[33923];
                
                r_data[33925] <= r_data[33924];
                
                r_data[33926] <= r_data[33925];
                
                r_data[33927] <= r_data[33926];
                
                r_data[33928] <= r_data[33927];
                
                r_data[33929] <= r_data[33928];
                
                r_data[33930] <= r_data[33929];
                
                r_data[33931] <= r_data[33930];
                
                r_data[33932] <= r_data[33931];
                
                r_data[33933] <= r_data[33932];
                
                r_data[33934] <= r_data[33933];
                
                r_data[33935] <= r_data[33934];
                
                r_data[33936] <= r_data[33935];
                
                r_data[33937] <= r_data[33936];
                
                r_data[33938] <= r_data[33937];
                
                r_data[33939] <= r_data[33938];
                
                r_data[33940] <= r_data[33939];
                
                r_data[33941] <= r_data[33940];
                
                r_data[33942] <= r_data[33941];
                
                r_data[33943] <= r_data[33942];
                
                r_data[33944] <= r_data[33943];
                
                r_data[33945] <= r_data[33944];
                
                r_data[33946] <= r_data[33945];
                
                r_data[33947] <= r_data[33946];
                
                r_data[33948] <= r_data[33947];
                
                r_data[33949] <= r_data[33948];
                
                r_data[33950] <= r_data[33949];
                
                r_data[33951] <= r_data[33950];
                
                r_data[33952] <= r_data[33951];
                
                r_data[33953] <= r_data[33952];
                
                r_data[33954] <= r_data[33953];
                
                r_data[33955] <= r_data[33954];
                
                r_data[33956] <= r_data[33955];
                
                r_data[33957] <= r_data[33956];
                
                r_data[33958] <= r_data[33957];
                
                r_data[33959] <= r_data[33958];
                
                r_data[33960] <= r_data[33959];
                
                r_data[33961] <= r_data[33960];
                
                r_data[33962] <= r_data[33961];
                
                r_data[33963] <= r_data[33962];
                
                r_data[33964] <= r_data[33963];
                
                r_data[33965] <= r_data[33964];
                
                r_data[33966] <= r_data[33965];
                
                r_data[33967] <= r_data[33966];
                
                r_data[33968] <= r_data[33967];
                
                r_data[33969] <= r_data[33968];
                
                r_data[33970] <= r_data[33969];
                
                r_data[33971] <= r_data[33970];
                
                r_data[33972] <= r_data[33971];
                
                r_data[33973] <= r_data[33972];
                
                r_data[33974] <= r_data[33973];
                
                r_data[33975] <= r_data[33974];
                
                r_data[33976] <= r_data[33975];
                
                r_data[33977] <= r_data[33976];
                
                r_data[33978] <= r_data[33977];
                
                r_data[33979] <= r_data[33978];
                
                r_data[33980] <= r_data[33979];
                
                r_data[33981] <= r_data[33980];
                
                r_data[33982] <= r_data[33981];
                
                r_data[33983] <= r_data[33982];
                
                r_data[33984] <= r_data[33983];
                
                r_data[33985] <= r_data[33984];
                
                r_data[33986] <= r_data[33985];
                
                r_data[33987] <= r_data[33986];
                
                r_data[33988] <= r_data[33987];
                
                r_data[33989] <= r_data[33988];
                
                r_data[33990] <= r_data[33989];
                
                r_data[33991] <= r_data[33990];
                
                r_data[33992] <= r_data[33991];
                
                r_data[33993] <= r_data[33992];
                
                r_data[33994] <= r_data[33993];
                
                r_data[33995] <= r_data[33994];
                
                r_data[33996] <= r_data[33995];
                
                r_data[33997] <= r_data[33996];
                
                r_data[33998] <= r_data[33997];
                
                r_data[33999] <= r_data[33998];
                
                r_data[34000] <= r_data[33999];
                
                r_data[34001] <= r_data[34000];
                
                r_data[34002] <= r_data[34001];
                
                r_data[34003] <= r_data[34002];
                
                r_data[34004] <= r_data[34003];
                
                r_data[34005] <= r_data[34004];
                
                r_data[34006] <= r_data[34005];
                
                r_data[34007] <= r_data[34006];
                
                r_data[34008] <= r_data[34007];
                
                r_data[34009] <= r_data[34008];
                
                r_data[34010] <= r_data[34009];
                
                r_data[34011] <= r_data[34010];
                
                r_data[34012] <= r_data[34011];
                
                r_data[34013] <= r_data[34012];
                
                r_data[34014] <= r_data[34013];
                
                r_data[34015] <= r_data[34014];
                
                r_data[34016] <= r_data[34015];
                
                r_data[34017] <= r_data[34016];
                
                r_data[34018] <= r_data[34017];
                
                r_data[34019] <= r_data[34018];
                
                r_data[34020] <= r_data[34019];
                
                r_data[34021] <= r_data[34020];
                
                r_data[34022] <= r_data[34021];
                
                r_data[34023] <= r_data[34022];
                
                r_data[34024] <= r_data[34023];
                
                r_data[34025] <= r_data[34024];
                
                r_data[34026] <= r_data[34025];
                
                r_data[34027] <= r_data[34026];
                
                r_data[34028] <= r_data[34027];
                
                r_data[34029] <= r_data[34028];
                
                r_data[34030] <= r_data[34029];
                
                r_data[34031] <= r_data[34030];
                
                r_data[34032] <= r_data[34031];
                
                r_data[34033] <= r_data[34032];
                
                r_data[34034] <= r_data[34033];
                
                r_data[34035] <= r_data[34034];
                
                r_data[34036] <= r_data[34035];
                
                r_data[34037] <= r_data[34036];
                
                r_data[34038] <= r_data[34037];
                
                r_data[34039] <= r_data[34038];
                
                r_data[34040] <= r_data[34039];
                
                r_data[34041] <= r_data[34040];
                
                r_data[34042] <= r_data[34041];
                
                r_data[34043] <= r_data[34042];
                
                r_data[34044] <= r_data[34043];
                
                r_data[34045] <= r_data[34044];
                
                r_data[34046] <= r_data[34045];
                
                r_data[34047] <= r_data[34046];
                
                r_data[34048] <= r_data[34047];
                
                r_data[34049] <= r_data[34048];
                
                r_data[34050] <= r_data[34049];
                
                r_data[34051] <= r_data[34050];
                
                r_data[34052] <= r_data[34051];
                
                r_data[34053] <= r_data[34052];
                
                r_data[34054] <= r_data[34053];
                
                r_data[34055] <= r_data[34054];
                
                r_data[34056] <= r_data[34055];
                
                r_data[34057] <= r_data[34056];
                
                r_data[34058] <= r_data[34057];
                
                r_data[34059] <= r_data[34058];
                
                r_data[34060] <= r_data[34059];
                
                r_data[34061] <= r_data[34060];
                
                r_data[34062] <= r_data[34061];
                
                r_data[34063] <= r_data[34062];
                
                r_data[34064] <= r_data[34063];
                
                r_data[34065] <= r_data[34064];
                
                r_data[34066] <= r_data[34065];
                
                r_data[34067] <= r_data[34066];
                
                r_data[34068] <= r_data[34067];
                
                r_data[34069] <= r_data[34068];
                
                r_data[34070] <= r_data[34069];
                
                r_data[34071] <= r_data[34070];
                
                r_data[34072] <= r_data[34071];
                
                r_data[34073] <= r_data[34072];
                
                r_data[34074] <= r_data[34073];
                
                r_data[34075] <= r_data[34074];
                
                r_data[34076] <= r_data[34075];
                
                r_data[34077] <= r_data[34076];
                
                r_data[34078] <= r_data[34077];
                
                r_data[34079] <= r_data[34078];
                
                r_data[34080] <= r_data[34079];
                
                r_data[34081] <= r_data[34080];
                
                r_data[34082] <= r_data[34081];
                
                r_data[34083] <= r_data[34082];
                
                r_data[34084] <= r_data[34083];
                
                r_data[34085] <= r_data[34084];
                
                r_data[34086] <= r_data[34085];
                
                r_data[34087] <= r_data[34086];
                
                r_data[34088] <= r_data[34087];
                
                r_data[34089] <= r_data[34088];
                
                r_data[34090] <= r_data[34089];
                
                r_data[34091] <= r_data[34090];
                
                r_data[34092] <= r_data[34091];
                
                r_data[34093] <= r_data[34092];
                
                r_data[34094] <= r_data[34093];
                
                r_data[34095] <= r_data[34094];
                
                r_data[34096] <= r_data[34095];
                
                r_data[34097] <= r_data[34096];
                
                r_data[34098] <= r_data[34097];
                
                r_data[34099] <= r_data[34098];
                
                r_data[34100] <= r_data[34099];
                
                r_data[34101] <= r_data[34100];
                
                r_data[34102] <= r_data[34101];
                
                r_data[34103] <= r_data[34102];
                
                r_data[34104] <= r_data[34103];
                
                r_data[34105] <= r_data[34104];
                
                r_data[34106] <= r_data[34105];
                
                r_data[34107] <= r_data[34106];
                
                r_data[34108] <= r_data[34107];
                
                r_data[34109] <= r_data[34108];
                
                r_data[34110] <= r_data[34109];
                
                r_data[34111] <= r_data[34110];
                
                r_data[34112] <= r_data[34111];
                
                r_data[34113] <= r_data[34112];
                
                r_data[34114] <= r_data[34113];
                
                r_data[34115] <= r_data[34114];
                
                r_data[34116] <= r_data[34115];
                
                r_data[34117] <= r_data[34116];
                
                r_data[34118] <= r_data[34117];
                
                r_data[34119] <= r_data[34118];
                
                r_data[34120] <= r_data[34119];
                
                r_data[34121] <= r_data[34120];
                
                r_data[34122] <= r_data[34121];
                
                r_data[34123] <= r_data[34122];
                
                r_data[34124] <= r_data[34123];
                
                r_data[34125] <= r_data[34124];
                
                r_data[34126] <= r_data[34125];
                
                r_data[34127] <= r_data[34126];
                
                r_data[34128] <= r_data[34127];
                
                r_data[34129] <= r_data[34128];
                
                r_data[34130] <= r_data[34129];
                
                r_data[34131] <= r_data[34130];
                
                r_data[34132] <= r_data[34131];
                
                r_data[34133] <= r_data[34132];
                
                r_data[34134] <= r_data[34133];
                
                r_data[34135] <= r_data[34134];
                
                r_data[34136] <= r_data[34135];
                
                r_data[34137] <= r_data[34136];
                
                r_data[34138] <= r_data[34137];
                
                r_data[34139] <= r_data[34138];
                
                r_data[34140] <= r_data[34139];
                
                r_data[34141] <= r_data[34140];
                
                r_data[34142] <= r_data[34141];
                
                r_data[34143] <= r_data[34142];
                
                r_data[34144] <= r_data[34143];
                
                r_data[34145] <= r_data[34144];
                
                r_data[34146] <= r_data[34145];
                
                r_data[34147] <= r_data[34146];
                
                r_data[34148] <= r_data[34147];
                
                r_data[34149] <= r_data[34148];
                
                r_data[34150] <= r_data[34149];
                
                r_data[34151] <= r_data[34150];
                
                r_data[34152] <= r_data[34151];
                
                r_data[34153] <= r_data[34152];
                
                r_data[34154] <= r_data[34153];
                
                r_data[34155] <= r_data[34154];
                
                r_data[34156] <= r_data[34155];
                
                r_data[34157] <= r_data[34156];
                
                r_data[34158] <= r_data[34157];
                
                r_data[34159] <= r_data[34158];
                
                r_data[34160] <= r_data[34159];
                
                r_data[34161] <= r_data[34160];
                
                r_data[34162] <= r_data[34161];
                
                r_data[34163] <= r_data[34162];
                
                r_data[34164] <= r_data[34163];
                
                r_data[34165] <= r_data[34164];
                
                r_data[34166] <= r_data[34165];
                
                r_data[34167] <= r_data[34166];
                
                r_data[34168] <= r_data[34167];
                
                r_data[34169] <= r_data[34168];
                
                r_data[34170] <= r_data[34169];
                
                r_data[34171] <= r_data[34170];
                
                r_data[34172] <= r_data[34171];
                
                r_data[34173] <= r_data[34172];
                
                r_data[34174] <= r_data[34173];
                
                r_data[34175] <= r_data[34174];
                
                r_data[34176] <= r_data[34175];
                
                r_data[34177] <= r_data[34176];
                
                r_data[34178] <= r_data[34177];
                
                r_data[34179] <= r_data[34178];
                
                r_data[34180] <= r_data[34179];
                
                r_data[34181] <= r_data[34180];
                
                r_data[34182] <= r_data[34181];
                
                r_data[34183] <= r_data[34182];
                
                r_data[34184] <= r_data[34183];
                
                r_data[34185] <= r_data[34184];
                
                r_data[34186] <= r_data[34185];
                
                r_data[34187] <= r_data[34186];
                
                r_data[34188] <= r_data[34187];
                
                r_data[34189] <= r_data[34188];
                
                r_data[34190] <= r_data[34189];
                
                r_data[34191] <= r_data[34190];
                
                r_data[34192] <= r_data[34191];
                
                r_data[34193] <= r_data[34192];
                
                r_data[34194] <= r_data[34193];
                
                r_data[34195] <= r_data[34194];
                
                r_data[34196] <= r_data[34195];
                
                r_data[34197] <= r_data[34196];
                
                r_data[34198] <= r_data[34197];
                
                r_data[34199] <= r_data[34198];
                
                r_data[34200] <= r_data[34199];
                
                r_data[34201] <= r_data[34200];
                
                r_data[34202] <= r_data[34201];
                
                r_data[34203] <= r_data[34202];
                
                r_data[34204] <= r_data[34203];
                
                r_data[34205] <= r_data[34204];
                
                r_data[34206] <= r_data[34205];
                
                r_data[34207] <= r_data[34206];
                
                r_data[34208] <= r_data[34207];
                
                r_data[34209] <= r_data[34208];
                
                r_data[34210] <= r_data[34209];
                
                r_data[34211] <= r_data[34210];
                
                r_data[34212] <= r_data[34211];
                
                r_data[34213] <= r_data[34212];
                
                r_data[34214] <= r_data[34213];
                
                r_data[34215] <= r_data[34214];
                
                r_data[34216] <= r_data[34215];
                
                r_data[34217] <= r_data[34216];
                
                r_data[34218] <= r_data[34217];
                
                r_data[34219] <= r_data[34218];
                
                r_data[34220] <= r_data[34219];
                
                r_data[34221] <= r_data[34220];
                
                r_data[34222] <= r_data[34221];
                
                r_data[34223] <= r_data[34222];
                
                r_data[34224] <= r_data[34223];
                
                r_data[34225] <= r_data[34224];
                
                r_data[34226] <= r_data[34225];
                
                r_data[34227] <= r_data[34226];
                
                r_data[34228] <= r_data[34227];
                
                r_data[34229] <= r_data[34228];
                
                r_data[34230] <= r_data[34229];
                
                r_data[34231] <= r_data[34230];
                
                r_data[34232] <= r_data[34231];
                
                r_data[34233] <= r_data[34232];
                
                r_data[34234] <= r_data[34233];
                
                r_data[34235] <= r_data[34234];
                
                r_data[34236] <= r_data[34235];
                
                r_data[34237] <= r_data[34236];
                
                r_data[34238] <= r_data[34237];
                
                r_data[34239] <= r_data[34238];
                
                r_data[34240] <= r_data[34239];
                
                r_data[34241] <= r_data[34240];
                
                r_data[34242] <= r_data[34241];
                
                r_data[34243] <= r_data[34242];
                
                r_data[34244] <= r_data[34243];
                
                r_data[34245] <= r_data[34244];
                
                r_data[34246] <= r_data[34245];
                
                r_data[34247] <= r_data[34246];
                
                r_data[34248] <= r_data[34247];
                
                r_data[34249] <= r_data[34248];
                
                r_data[34250] <= r_data[34249];
                
                r_data[34251] <= r_data[34250];
                
                r_data[34252] <= r_data[34251];
                
                r_data[34253] <= r_data[34252];
                
                r_data[34254] <= r_data[34253];
                
                r_data[34255] <= r_data[34254];
                
                r_data[34256] <= r_data[34255];
                
                r_data[34257] <= r_data[34256];
                
                r_data[34258] <= r_data[34257];
                
                r_data[34259] <= r_data[34258];
                
                r_data[34260] <= r_data[34259];
                
                r_data[34261] <= r_data[34260];
                
                r_data[34262] <= r_data[34261];
                
                r_data[34263] <= r_data[34262];
                
                r_data[34264] <= r_data[34263];
                
                r_data[34265] <= r_data[34264];
                
                r_data[34266] <= r_data[34265];
                
                r_data[34267] <= r_data[34266];
                
                r_data[34268] <= r_data[34267];
                
                r_data[34269] <= r_data[34268];
                
                r_data[34270] <= r_data[34269];
                
                r_data[34271] <= r_data[34270];
                
                r_data[34272] <= r_data[34271];
                
                r_data[34273] <= r_data[34272];
                
                r_data[34274] <= r_data[34273];
                
                r_data[34275] <= r_data[34274];
                
                r_data[34276] <= r_data[34275];
                
                r_data[34277] <= r_data[34276];
                
                r_data[34278] <= r_data[34277];
                
                r_data[34279] <= r_data[34278];
                
                r_data[34280] <= r_data[34279];
                
                r_data[34281] <= r_data[34280];
                
                r_data[34282] <= r_data[34281];
                
                r_data[34283] <= r_data[34282];
                
                r_data[34284] <= r_data[34283];
                
                r_data[34285] <= r_data[34284];
                
                r_data[34286] <= r_data[34285];
                
                r_data[34287] <= r_data[34286];
                
                r_data[34288] <= r_data[34287];
                
                r_data[34289] <= r_data[34288];
                
                r_data[34290] <= r_data[34289];
                
                r_data[34291] <= r_data[34290];
                
                r_data[34292] <= r_data[34291];
                
                r_data[34293] <= r_data[34292];
                
                r_data[34294] <= r_data[34293];
                
                r_data[34295] <= r_data[34294];
                
                r_data[34296] <= r_data[34295];
                
                r_data[34297] <= r_data[34296];
                
                r_data[34298] <= r_data[34297];
                
                r_data[34299] <= r_data[34298];
                
                r_data[34300] <= r_data[34299];
                
                r_data[34301] <= r_data[34300];
                
                r_data[34302] <= r_data[34301];
                
                r_data[34303] <= r_data[34302];
                
                r_data[34304] <= r_data[34303];
                
                r_data[34305] <= r_data[34304];
                
                r_data[34306] <= r_data[34305];
                
                r_data[34307] <= r_data[34306];
                
                r_data[34308] <= r_data[34307];
                
                r_data[34309] <= r_data[34308];
                
                r_data[34310] <= r_data[34309];
                
                r_data[34311] <= r_data[34310];
                
                r_data[34312] <= r_data[34311];
                
                r_data[34313] <= r_data[34312];
                
                r_data[34314] <= r_data[34313];
                
                r_data[34315] <= r_data[34314];
                
                r_data[34316] <= r_data[34315];
                
                r_data[34317] <= r_data[34316];
                
                r_data[34318] <= r_data[34317];
                
                r_data[34319] <= r_data[34318];
                
                r_data[34320] <= r_data[34319];
                
                r_data[34321] <= r_data[34320];
                
                r_data[34322] <= r_data[34321];
                
                r_data[34323] <= r_data[34322];
                
                r_data[34324] <= r_data[34323];
                
                r_data[34325] <= r_data[34324];
                
                r_data[34326] <= r_data[34325];
                
                r_data[34327] <= r_data[34326];
                
                r_data[34328] <= r_data[34327];
                
                r_data[34329] <= r_data[34328];
                
                r_data[34330] <= r_data[34329];
                
                r_data[34331] <= r_data[34330];
                
                r_data[34332] <= r_data[34331];
                
                r_data[34333] <= r_data[34332];
                
                r_data[34334] <= r_data[34333];
                
                r_data[34335] <= r_data[34334];
                
                r_data[34336] <= r_data[34335];
                
                r_data[34337] <= r_data[34336];
                
                r_data[34338] <= r_data[34337];
                
                r_data[34339] <= r_data[34338];
                
                r_data[34340] <= r_data[34339];
                
                r_data[34341] <= r_data[34340];
                
                r_data[34342] <= r_data[34341];
                
                r_data[34343] <= r_data[34342];
                
                r_data[34344] <= r_data[34343];
                
                r_data[34345] <= r_data[34344];
                
                r_data[34346] <= r_data[34345];
                
                r_data[34347] <= r_data[34346];
                
                r_data[34348] <= r_data[34347];
                
                r_data[34349] <= r_data[34348];
                
                r_data[34350] <= r_data[34349];
                
                r_data[34351] <= r_data[34350];
                
                r_data[34352] <= r_data[34351];
                
                r_data[34353] <= r_data[34352];
                
                r_data[34354] <= r_data[34353];
                
                r_data[34355] <= r_data[34354];
                
                r_data[34356] <= r_data[34355];
                
                r_data[34357] <= r_data[34356];
                
                r_data[34358] <= r_data[34357];
                
                r_data[34359] <= r_data[34358];
                
                r_data[34360] <= r_data[34359];
                
                r_data[34361] <= r_data[34360];
                
                r_data[34362] <= r_data[34361];
                
                r_data[34363] <= r_data[34362];
                
                r_data[34364] <= r_data[34363];
                
                r_data[34365] <= r_data[34364];
                
                r_data[34366] <= r_data[34365];
                
                r_data[34367] <= r_data[34366];
                
                r_data[34368] <= r_data[34367];
                
                r_data[34369] <= r_data[34368];
                
                r_data[34370] <= r_data[34369];
                
                r_data[34371] <= r_data[34370];
                
                r_data[34372] <= r_data[34371];
                
                r_data[34373] <= r_data[34372];
                
                r_data[34374] <= r_data[34373];
                
                r_data[34375] <= r_data[34374];
                
                r_data[34376] <= r_data[34375];
                
                r_data[34377] <= r_data[34376];
                
                r_data[34378] <= r_data[34377];
                
                r_data[34379] <= r_data[34378];
                
                r_data[34380] <= r_data[34379];
                
                r_data[34381] <= r_data[34380];
                
                r_data[34382] <= r_data[34381];
                
                r_data[34383] <= r_data[34382];
                
                r_data[34384] <= r_data[34383];
                
                r_data[34385] <= r_data[34384];
                
                r_data[34386] <= r_data[34385];
                
                r_data[34387] <= r_data[34386];
                
                r_data[34388] <= r_data[34387];
                
                r_data[34389] <= r_data[34388];
                
                r_data[34390] <= r_data[34389];
                
                r_data[34391] <= r_data[34390];
                
                r_data[34392] <= r_data[34391];
                
                r_data[34393] <= r_data[34392];
                
                r_data[34394] <= r_data[34393];
                
                r_data[34395] <= r_data[34394];
                
                r_data[34396] <= r_data[34395];
                
                r_data[34397] <= r_data[34396];
                
                r_data[34398] <= r_data[34397];
                
                r_data[34399] <= r_data[34398];
                
                r_data[34400] <= r_data[34399];
                
                r_data[34401] <= r_data[34400];
                
                r_data[34402] <= r_data[34401];
                
                r_data[34403] <= r_data[34402];
                
                r_data[34404] <= r_data[34403];
                
                r_data[34405] <= r_data[34404];
                
                r_data[34406] <= r_data[34405];
                
                r_data[34407] <= r_data[34406];
                
                r_data[34408] <= r_data[34407];
                
                r_data[34409] <= r_data[34408];
                
                r_data[34410] <= r_data[34409];
                
                r_data[34411] <= r_data[34410];
                
                r_data[34412] <= r_data[34411];
                
                r_data[34413] <= r_data[34412];
                
                r_data[34414] <= r_data[34413];
                
                r_data[34415] <= r_data[34414];
                
                r_data[34416] <= r_data[34415];
                
                r_data[34417] <= r_data[34416];
                
                r_data[34418] <= r_data[34417];
                
                r_data[34419] <= r_data[34418];
                
                r_data[34420] <= r_data[34419];
                
                r_data[34421] <= r_data[34420];
                
                r_data[34422] <= r_data[34421];
                
                r_data[34423] <= r_data[34422];
                
                r_data[34424] <= r_data[34423];
                
                r_data[34425] <= r_data[34424];
                
                r_data[34426] <= r_data[34425];
                
                r_data[34427] <= r_data[34426];
                
                r_data[34428] <= r_data[34427];
                
                r_data[34429] <= r_data[34428];
                
                r_data[34430] <= r_data[34429];
                
                r_data[34431] <= r_data[34430];
                
                r_data[34432] <= r_data[34431];
                
                r_data[34433] <= r_data[34432];
                
                r_data[34434] <= r_data[34433];
                
                r_data[34435] <= r_data[34434];
                
                r_data[34436] <= r_data[34435];
                
                r_data[34437] <= r_data[34436];
                
                r_data[34438] <= r_data[34437];
                
                r_data[34439] <= r_data[34438];
                
                r_data[34440] <= r_data[34439];
                
                r_data[34441] <= r_data[34440];
                
                r_data[34442] <= r_data[34441];
                
                r_data[34443] <= r_data[34442];
                
                r_data[34444] <= r_data[34443];
                
                r_data[34445] <= r_data[34444];
                
                r_data[34446] <= r_data[34445];
                
                r_data[34447] <= r_data[34446];
                
                r_data[34448] <= r_data[34447];
                
                r_data[34449] <= r_data[34448];
                
                r_data[34450] <= r_data[34449];
                
                r_data[34451] <= r_data[34450];
                
                r_data[34452] <= r_data[34451];
                
                r_data[34453] <= r_data[34452];
                
                r_data[34454] <= r_data[34453];
                
                r_data[34455] <= r_data[34454];
                
                r_data[34456] <= r_data[34455];
                
                r_data[34457] <= r_data[34456];
                
                r_data[34458] <= r_data[34457];
                
                r_data[34459] <= r_data[34458];
                
                r_data[34460] <= r_data[34459];
                
                r_data[34461] <= r_data[34460];
                
                r_data[34462] <= r_data[34461];
                
                r_data[34463] <= r_data[34462];
                
                r_data[34464] <= r_data[34463];
                
                r_data[34465] <= r_data[34464];
                
                r_data[34466] <= r_data[34465];
                
                r_data[34467] <= r_data[34466];
                
                r_data[34468] <= r_data[34467];
                
                r_data[34469] <= r_data[34468];
                
                r_data[34470] <= r_data[34469];
                
                r_data[34471] <= r_data[34470];
                
                r_data[34472] <= r_data[34471];
                
                r_data[34473] <= r_data[34472];
                
                r_data[34474] <= r_data[34473];
                
                r_data[34475] <= r_data[34474];
                
                r_data[34476] <= r_data[34475];
                
                r_data[34477] <= r_data[34476];
                
                r_data[34478] <= r_data[34477];
                
                r_data[34479] <= r_data[34478];
                
                r_data[34480] <= r_data[34479];
                
                r_data[34481] <= r_data[34480];
                
                r_data[34482] <= r_data[34481];
                
                r_data[34483] <= r_data[34482];
                
                r_data[34484] <= r_data[34483];
                
                r_data[34485] <= r_data[34484];
                
                r_data[34486] <= r_data[34485];
                
                r_data[34487] <= r_data[34486];
                
                r_data[34488] <= r_data[34487];
                
                r_data[34489] <= r_data[34488];
                
                r_data[34490] <= r_data[34489];
                
                r_data[34491] <= r_data[34490];
                
                r_data[34492] <= r_data[34491];
                
                r_data[34493] <= r_data[34492];
                
                r_data[34494] <= r_data[34493];
                
                r_data[34495] <= r_data[34494];
                
                r_data[34496] <= r_data[34495];
                
                r_data[34497] <= r_data[34496];
                
                r_data[34498] <= r_data[34497];
                
                r_data[34499] <= r_data[34498];
                
                r_data[34500] <= r_data[34499];
                
                r_data[34501] <= r_data[34500];
                
                r_data[34502] <= r_data[34501];
                
                r_data[34503] <= r_data[34502];
                
                r_data[34504] <= r_data[34503];
                
                r_data[34505] <= r_data[34504];
                
                r_data[34506] <= r_data[34505];
                
                r_data[34507] <= r_data[34506];
                
                r_data[34508] <= r_data[34507];
                
                r_data[34509] <= r_data[34508];
                
                r_data[34510] <= r_data[34509];
                
                r_data[34511] <= r_data[34510];
                
                r_data[34512] <= r_data[34511];
                
                r_data[34513] <= r_data[34512];
                
                r_data[34514] <= r_data[34513];
                
                r_data[34515] <= r_data[34514];
                
                r_data[34516] <= r_data[34515];
                
                r_data[34517] <= r_data[34516];
                
                r_data[34518] <= r_data[34517];
                
                r_data[34519] <= r_data[34518];
                
                r_data[34520] <= r_data[34519];
                
                r_data[34521] <= r_data[34520];
                
                r_data[34522] <= r_data[34521];
                
                r_data[34523] <= r_data[34522];
                
                r_data[34524] <= r_data[34523];
                
                r_data[34525] <= r_data[34524];
                
                r_data[34526] <= r_data[34525];
                
                r_data[34527] <= r_data[34526];
                
                r_data[34528] <= r_data[34527];
                
                r_data[34529] <= r_data[34528];
                
                r_data[34530] <= r_data[34529];
                
                r_data[34531] <= r_data[34530];
                
                r_data[34532] <= r_data[34531];
                
                r_data[34533] <= r_data[34532];
                
                r_data[34534] <= r_data[34533];
                
                r_data[34535] <= r_data[34534];
                
                r_data[34536] <= r_data[34535];
                
                r_data[34537] <= r_data[34536];
                
                r_data[34538] <= r_data[34537];
                
                r_data[34539] <= r_data[34538];
                
                r_data[34540] <= r_data[34539];
                
                r_data[34541] <= r_data[34540];
                
                r_data[34542] <= r_data[34541];
                
                r_data[34543] <= r_data[34542];
                
                r_data[34544] <= r_data[34543];
                
                r_data[34545] <= r_data[34544];
                
                r_data[34546] <= r_data[34545];
                
                r_data[34547] <= r_data[34546];
                
                r_data[34548] <= r_data[34547];
                
                r_data[34549] <= r_data[34548];
                
                r_data[34550] <= r_data[34549];
                
                r_data[34551] <= r_data[34550];
                
                r_data[34552] <= r_data[34551];
                
                r_data[34553] <= r_data[34552];
                
                r_data[34554] <= r_data[34553];
                
                r_data[34555] <= r_data[34554];
                
                r_data[34556] <= r_data[34555];
                
                r_data[34557] <= r_data[34556];
                
                r_data[34558] <= r_data[34557];
                
                r_data[34559] <= r_data[34558];
                
                r_data[34560] <= r_data[34559];
                
                r_data[34561] <= r_data[34560];
                
                r_data[34562] <= r_data[34561];
                
                r_data[34563] <= r_data[34562];
                
                r_data[34564] <= r_data[34563];
                
                r_data[34565] <= r_data[34564];
                
                r_data[34566] <= r_data[34565];
                
                r_data[34567] <= r_data[34566];
                
                r_data[34568] <= r_data[34567];
                
                r_data[34569] <= r_data[34568];
                
                r_data[34570] <= r_data[34569];
                
                r_data[34571] <= r_data[34570];
                
                r_data[34572] <= r_data[34571];
                
                r_data[34573] <= r_data[34572];
                
                r_data[34574] <= r_data[34573];
                
                r_data[34575] <= r_data[34574];
                
                r_data[34576] <= r_data[34575];
                
                r_data[34577] <= r_data[34576];
                
                r_data[34578] <= r_data[34577];
                
                r_data[34579] <= r_data[34578];
                
                r_data[34580] <= r_data[34579];
                
                r_data[34581] <= r_data[34580];
                
                r_data[34582] <= r_data[34581];
                
                r_data[34583] <= r_data[34582];
                
                r_data[34584] <= r_data[34583];
                
                r_data[34585] <= r_data[34584];
                
                r_data[34586] <= r_data[34585];
                
                r_data[34587] <= r_data[34586];
                
                r_data[34588] <= r_data[34587];
                
                r_data[34589] <= r_data[34588];
                
                r_data[34590] <= r_data[34589];
                
                r_data[34591] <= r_data[34590];
                
                r_data[34592] <= r_data[34591];
                
                r_data[34593] <= r_data[34592];
                
                r_data[34594] <= r_data[34593];
                
                r_data[34595] <= r_data[34594];
                
                r_data[34596] <= r_data[34595];
                
                r_data[34597] <= r_data[34596];
                
                r_data[34598] <= r_data[34597];
                
                r_data[34599] <= r_data[34598];
                
                r_data[34600] <= r_data[34599];
                
                r_data[34601] <= r_data[34600];
                
                r_data[34602] <= r_data[34601];
                
                r_data[34603] <= r_data[34602];
                
                r_data[34604] <= r_data[34603];
                
                r_data[34605] <= r_data[34604];
                
                r_data[34606] <= r_data[34605];
                
                r_data[34607] <= r_data[34606];
                
                r_data[34608] <= r_data[34607];
                
                r_data[34609] <= r_data[34608];
                
                r_data[34610] <= r_data[34609];
                
                r_data[34611] <= r_data[34610];
                
                r_data[34612] <= r_data[34611];
                
                r_data[34613] <= r_data[34612];
                
                r_data[34614] <= r_data[34613];
                
                r_data[34615] <= r_data[34614];
                
                r_data[34616] <= r_data[34615];
                
                r_data[34617] <= r_data[34616];
                
                r_data[34618] <= r_data[34617];
                
                r_data[34619] <= r_data[34618];
                
                r_data[34620] <= r_data[34619];
                
                r_data[34621] <= r_data[34620];
                
                r_data[34622] <= r_data[34621];
                
                r_data[34623] <= r_data[34622];
                
                r_data[34624] <= r_data[34623];
                
                r_data[34625] <= r_data[34624];
                
                r_data[34626] <= r_data[34625];
                
                r_data[34627] <= r_data[34626];
                
                r_data[34628] <= r_data[34627];
                
                r_data[34629] <= r_data[34628];
                
                r_data[34630] <= r_data[34629];
                
                r_data[34631] <= r_data[34630];
                
                r_data[34632] <= r_data[34631];
                
                r_data[34633] <= r_data[34632];
                
                r_data[34634] <= r_data[34633];
                
                r_data[34635] <= r_data[34634];
                
                r_data[34636] <= r_data[34635];
                
                r_data[34637] <= r_data[34636];
                
                r_data[34638] <= r_data[34637];
                
                r_data[34639] <= r_data[34638];
                
                r_data[34640] <= r_data[34639];
                
                r_data[34641] <= r_data[34640];
                
                r_data[34642] <= r_data[34641];
                
                r_data[34643] <= r_data[34642];
                
                r_data[34644] <= r_data[34643];
                
                r_data[34645] <= r_data[34644];
                
                r_data[34646] <= r_data[34645];
                
                r_data[34647] <= r_data[34646];
                
                r_data[34648] <= r_data[34647];
                
                r_data[34649] <= r_data[34648];
                
                r_data[34650] <= r_data[34649];
                
                r_data[34651] <= r_data[34650];
                
                r_data[34652] <= r_data[34651];
                
                r_data[34653] <= r_data[34652];
                
                r_data[34654] <= r_data[34653];
                
                r_data[34655] <= r_data[34654];
                
                r_data[34656] <= r_data[34655];
                
                r_data[34657] <= r_data[34656];
                
                r_data[34658] <= r_data[34657];
                
                r_data[34659] <= r_data[34658];
                
                r_data[34660] <= r_data[34659];
                
                r_data[34661] <= r_data[34660];
                
                r_data[34662] <= r_data[34661];
                
                r_data[34663] <= r_data[34662];
                
                r_data[34664] <= r_data[34663];
                
                r_data[34665] <= r_data[34664];
                
                r_data[34666] <= r_data[34665];
                
                r_data[34667] <= r_data[34666];
                
                r_data[34668] <= r_data[34667];
                
                r_data[34669] <= r_data[34668];
                
                r_data[34670] <= r_data[34669];
                
                r_data[34671] <= r_data[34670];
                
                r_data[34672] <= r_data[34671];
                
                r_data[34673] <= r_data[34672];
                
                r_data[34674] <= r_data[34673];
                
                r_data[34675] <= r_data[34674];
                
                r_data[34676] <= r_data[34675];
                
                r_data[34677] <= r_data[34676];
                
                r_data[34678] <= r_data[34677];
                
                r_data[34679] <= r_data[34678];
                
                r_data[34680] <= r_data[34679];
                
                r_data[34681] <= r_data[34680];
                
                r_data[34682] <= r_data[34681];
                
                r_data[34683] <= r_data[34682];
                
                r_data[34684] <= r_data[34683];
                
                r_data[34685] <= r_data[34684];
                
                r_data[34686] <= r_data[34685];
                
                r_data[34687] <= r_data[34686];
                
                r_data[34688] <= r_data[34687];
                
                r_data[34689] <= r_data[34688];
                
                r_data[34690] <= r_data[34689];
                
                r_data[34691] <= r_data[34690];
                
                r_data[34692] <= r_data[34691];
                
                r_data[34693] <= r_data[34692];
                
                r_data[34694] <= r_data[34693];
                
                r_data[34695] <= r_data[34694];
                
                r_data[34696] <= r_data[34695];
                
                r_data[34697] <= r_data[34696];
                
                r_data[34698] <= r_data[34697];
                
                r_data[34699] <= r_data[34698];
                
                r_data[34700] <= r_data[34699];
                
                r_data[34701] <= r_data[34700];
                
                r_data[34702] <= r_data[34701];
                
                r_data[34703] <= r_data[34702];
                
                r_data[34704] <= r_data[34703];
                
                r_data[34705] <= r_data[34704];
                
                r_data[34706] <= r_data[34705];
                
                r_data[34707] <= r_data[34706];
                
                r_data[34708] <= r_data[34707];
                
                r_data[34709] <= r_data[34708];
                
                r_data[34710] <= r_data[34709];
                
                r_data[34711] <= r_data[34710];
                
                r_data[34712] <= r_data[34711];
                
                r_data[34713] <= r_data[34712];
                
                r_data[34714] <= r_data[34713];
                
                r_data[34715] <= r_data[34714];
                
                r_data[34716] <= r_data[34715];
                
                r_data[34717] <= r_data[34716];
                
                r_data[34718] <= r_data[34717];
                
                r_data[34719] <= r_data[34718];
                
                r_data[34720] <= r_data[34719];
                
                r_data[34721] <= r_data[34720];
                
                r_data[34722] <= r_data[34721];
                
                r_data[34723] <= r_data[34722];
                
                r_data[34724] <= r_data[34723];
                
                r_data[34725] <= r_data[34724];
                
                r_data[34726] <= r_data[34725];
                
                r_data[34727] <= r_data[34726];
                
                r_data[34728] <= r_data[34727];
                
                r_data[34729] <= r_data[34728];
                
                r_data[34730] <= r_data[34729];
                
                r_data[34731] <= r_data[34730];
                
                r_data[34732] <= r_data[34731];
                
                r_data[34733] <= r_data[34732];
                
                r_data[34734] <= r_data[34733];
                
                r_data[34735] <= r_data[34734];
                
                r_data[34736] <= r_data[34735];
                
                r_data[34737] <= r_data[34736];
                
                r_data[34738] <= r_data[34737];
                
                r_data[34739] <= r_data[34738];
                
                r_data[34740] <= r_data[34739];
                
                r_data[34741] <= r_data[34740];
                
                r_data[34742] <= r_data[34741];
                
                r_data[34743] <= r_data[34742];
                
                r_data[34744] <= r_data[34743];
                
                r_data[34745] <= r_data[34744];
                
                r_data[34746] <= r_data[34745];
                
                r_data[34747] <= r_data[34746];
                
                r_data[34748] <= r_data[34747];
                
                r_data[34749] <= r_data[34748];
                
                r_data[34750] <= r_data[34749];
                
                r_data[34751] <= r_data[34750];
                
                r_data[34752] <= r_data[34751];
                
                r_data[34753] <= r_data[34752];
                
                r_data[34754] <= r_data[34753];
                
                r_data[34755] <= r_data[34754];
                
                r_data[34756] <= r_data[34755];
                
                r_data[34757] <= r_data[34756];
                
                r_data[34758] <= r_data[34757];
                
                r_data[34759] <= r_data[34758];
                
                r_data[34760] <= r_data[34759];
                
                r_data[34761] <= r_data[34760];
                
                r_data[34762] <= r_data[34761];
                
                r_data[34763] <= r_data[34762];
                
                r_data[34764] <= r_data[34763];
                
                r_data[34765] <= r_data[34764];
                
                r_data[34766] <= r_data[34765];
                
                r_data[34767] <= r_data[34766];
                
                r_data[34768] <= r_data[34767];
                
                r_data[34769] <= r_data[34768];
                
                r_data[34770] <= r_data[34769];
                
                r_data[34771] <= r_data[34770];
                
                r_data[34772] <= r_data[34771];
                
                r_data[34773] <= r_data[34772];
                
                r_data[34774] <= r_data[34773];
                
                r_data[34775] <= r_data[34774];
                
                r_data[34776] <= r_data[34775];
                
                r_data[34777] <= r_data[34776];
                
                r_data[34778] <= r_data[34777];
                
                r_data[34779] <= r_data[34778];
                
                r_data[34780] <= r_data[34779];
                
                r_data[34781] <= r_data[34780];
                
                r_data[34782] <= r_data[34781];
                
                r_data[34783] <= r_data[34782];
                
                r_data[34784] <= r_data[34783];
                
                r_data[34785] <= r_data[34784];
                
                r_data[34786] <= r_data[34785];
                
                r_data[34787] <= r_data[34786];
                
                r_data[34788] <= r_data[34787];
                
                r_data[34789] <= r_data[34788];
                
                r_data[34790] <= r_data[34789];
                
                r_data[34791] <= r_data[34790];
                
                r_data[34792] <= r_data[34791];
                
                r_data[34793] <= r_data[34792];
                
                r_data[34794] <= r_data[34793];
                
                r_data[34795] <= r_data[34794];
                
                r_data[34796] <= r_data[34795];
                
                r_data[34797] <= r_data[34796];
                
                r_data[34798] <= r_data[34797];
                
                r_data[34799] <= r_data[34798];
                
                r_data[34800] <= r_data[34799];
                
                r_data[34801] <= r_data[34800];
                
                r_data[34802] <= r_data[34801];
                
                r_data[34803] <= r_data[34802];
                
                r_data[34804] <= r_data[34803];
                
                r_data[34805] <= r_data[34804];
                
                r_data[34806] <= r_data[34805];
                
                r_data[34807] <= r_data[34806];
                
                r_data[34808] <= r_data[34807];
                
                r_data[34809] <= r_data[34808];
                
                r_data[34810] <= r_data[34809];
                
                r_data[34811] <= r_data[34810];
                
                r_data[34812] <= r_data[34811];
                
                r_data[34813] <= r_data[34812];
                
                r_data[34814] <= r_data[34813];
                
                r_data[34815] <= r_data[34814];
                
                r_data[34816] <= r_data[34815];
                
                r_data[34817] <= r_data[34816];
                
                r_data[34818] <= r_data[34817];
                
                r_data[34819] <= r_data[34818];
                
                r_data[34820] <= r_data[34819];
                
                r_data[34821] <= r_data[34820];
                
                r_data[34822] <= r_data[34821];
                
                r_data[34823] <= r_data[34822];
                
                r_data[34824] <= r_data[34823];
                
                r_data[34825] <= r_data[34824];
                
                r_data[34826] <= r_data[34825];
                
                r_data[34827] <= r_data[34826];
                
                r_data[34828] <= r_data[34827];
                
                r_data[34829] <= r_data[34828];
                
                r_data[34830] <= r_data[34829];
                
                r_data[34831] <= r_data[34830];
                
                r_data[34832] <= r_data[34831];
                
                r_data[34833] <= r_data[34832];
                
                r_data[34834] <= r_data[34833];
                
                r_data[34835] <= r_data[34834];
                
                r_data[34836] <= r_data[34835];
                
                r_data[34837] <= r_data[34836];
                
                r_data[34838] <= r_data[34837];
                
                r_data[34839] <= r_data[34838];
                
                r_data[34840] <= r_data[34839];
                
                r_data[34841] <= r_data[34840];
                
                r_data[34842] <= r_data[34841];
                
                r_data[34843] <= r_data[34842];
                
                r_data[34844] <= r_data[34843];
                
                r_data[34845] <= r_data[34844];
                
                r_data[34846] <= r_data[34845];
                
                r_data[34847] <= r_data[34846];
                
                r_data[34848] <= r_data[34847];
                
                r_data[34849] <= r_data[34848];
                
                r_data[34850] <= r_data[34849];
                
                r_data[34851] <= r_data[34850];
                
                r_data[34852] <= r_data[34851];
                
                r_data[34853] <= r_data[34852];
                
                r_data[34854] <= r_data[34853];
                
                r_data[34855] <= r_data[34854];
                
                r_data[34856] <= r_data[34855];
                
                r_data[34857] <= r_data[34856];
                
                r_data[34858] <= r_data[34857];
                
                r_data[34859] <= r_data[34858];
                
                r_data[34860] <= r_data[34859];
                
                r_data[34861] <= r_data[34860];
                
                r_data[34862] <= r_data[34861];
                
                r_data[34863] <= r_data[34862];
                
                r_data[34864] <= r_data[34863];
                
                r_data[34865] <= r_data[34864];
                
                r_data[34866] <= r_data[34865];
                
                r_data[34867] <= r_data[34866];
                
                r_data[34868] <= r_data[34867];
                
                r_data[34869] <= r_data[34868];
                
                r_data[34870] <= r_data[34869];
                
                r_data[34871] <= r_data[34870];
                
                r_data[34872] <= r_data[34871];
                
                r_data[34873] <= r_data[34872];
                
                r_data[34874] <= r_data[34873];
                
                r_data[34875] <= r_data[34874];
                
                r_data[34876] <= r_data[34875];
                
                r_data[34877] <= r_data[34876];
                
                r_data[34878] <= r_data[34877];
                
                r_data[34879] <= r_data[34878];
                
                r_data[34880] <= r_data[34879];
                
                r_data[34881] <= r_data[34880];
                
                r_data[34882] <= r_data[34881];
                
                r_data[34883] <= r_data[34882];
                
                r_data[34884] <= r_data[34883];
                
                r_data[34885] <= r_data[34884];
                
                r_data[34886] <= r_data[34885];
                
                r_data[34887] <= r_data[34886];
                
                r_data[34888] <= r_data[34887];
                
                r_data[34889] <= r_data[34888];
                
                r_data[34890] <= r_data[34889];
                
                r_data[34891] <= r_data[34890];
                
                r_data[34892] <= r_data[34891];
                
                r_data[34893] <= r_data[34892];
                
                r_data[34894] <= r_data[34893];
                
                r_data[34895] <= r_data[34894];
                
                r_data[34896] <= r_data[34895];
                
                r_data[34897] <= r_data[34896];
                
                r_data[34898] <= r_data[34897];
                
                r_data[34899] <= r_data[34898];
                
                r_data[34900] <= r_data[34899];
                
                r_data[34901] <= r_data[34900];
                
                r_data[34902] <= r_data[34901];
                
                r_data[34903] <= r_data[34902];
                
                r_data[34904] <= r_data[34903];
                
                r_data[34905] <= r_data[34904];
                
                r_data[34906] <= r_data[34905];
                
                r_data[34907] <= r_data[34906];
                
                r_data[34908] <= r_data[34907];
                
                r_data[34909] <= r_data[34908];
                
                r_data[34910] <= r_data[34909];
                
                r_data[34911] <= r_data[34910];
                
                r_data[34912] <= r_data[34911];
                
                r_data[34913] <= r_data[34912];
                
                r_data[34914] <= r_data[34913];
                
                r_data[34915] <= r_data[34914];
                
                r_data[34916] <= r_data[34915];
                
                r_data[34917] <= r_data[34916];
                
                r_data[34918] <= r_data[34917];
                
                r_data[34919] <= r_data[34918];
                
                r_data[34920] <= r_data[34919];
                
                r_data[34921] <= r_data[34920];
                
                r_data[34922] <= r_data[34921];
                
                r_data[34923] <= r_data[34922];
                
                r_data[34924] <= r_data[34923];
                
                r_data[34925] <= r_data[34924];
                
                r_data[34926] <= r_data[34925];
                
                r_data[34927] <= r_data[34926];
                
                r_data[34928] <= r_data[34927];
                
                r_data[34929] <= r_data[34928];
                
                r_data[34930] <= r_data[34929];
                
                r_data[34931] <= r_data[34930];
                
                r_data[34932] <= r_data[34931];
                
                r_data[34933] <= r_data[34932];
                
                r_data[34934] <= r_data[34933];
                
                r_data[34935] <= r_data[34934];
                
                r_data[34936] <= r_data[34935];
                
                r_data[34937] <= r_data[34936];
                
                r_data[34938] <= r_data[34937];
                
                r_data[34939] <= r_data[34938];
                
                r_data[34940] <= r_data[34939];
                
                r_data[34941] <= r_data[34940];
                
                r_data[34942] <= r_data[34941];
                
                r_data[34943] <= r_data[34942];
                
                r_data[34944] <= r_data[34943];
                
                r_data[34945] <= r_data[34944];
                
                r_data[34946] <= r_data[34945];
                
                r_data[34947] <= r_data[34946];
                
                r_data[34948] <= r_data[34947];
                
                r_data[34949] <= r_data[34948];
                
                r_data[34950] <= r_data[34949];
                
                r_data[34951] <= r_data[34950];
                
                r_data[34952] <= r_data[34951];
                
                r_data[34953] <= r_data[34952];
                
                r_data[34954] <= r_data[34953];
                
                r_data[34955] <= r_data[34954];
                
                r_data[34956] <= r_data[34955];
                
                r_data[34957] <= r_data[34956];
                
                r_data[34958] <= r_data[34957];
                
                r_data[34959] <= r_data[34958];
                
                r_data[34960] <= r_data[34959];
                
                r_data[34961] <= r_data[34960];
                
                r_data[34962] <= r_data[34961];
                
                r_data[34963] <= r_data[34962];
                
                r_data[34964] <= r_data[34963];
                
                r_data[34965] <= r_data[34964];
                
                r_data[34966] <= r_data[34965];
                
                r_data[34967] <= r_data[34966];
                
                r_data[34968] <= r_data[34967];
                
                r_data[34969] <= r_data[34968];
                
                r_data[34970] <= r_data[34969];
                
                r_data[34971] <= r_data[34970];
                
                r_data[34972] <= r_data[34971];
                
                r_data[34973] <= r_data[34972];
                
                r_data[34974] <= r_data[34973];
                
                r_data[34975] <= r_data[34974];
                
                r_data[34976] <= r_data[34975];
                
                r_data[34977] <= r_data[34976];
                
                r_data[34978] <= r_data[34977];
                
                r_data[34979] <= r_data[34978];
                
                r_data[34980] <= r_data[34979];
                
                r_data[34981] <= r_data[34980];
                
                r_data[34982] <= r_data[34981];
                
                r_data[34983] <= r_data[34982];
                
                r_data[34984] <= r_data[34983];
                
                r_data[34985] <= r_data[34984];
                
                r_data[34986] <= r_data[34985];
                
                r_data[34987] <= r_data[34986];
                
                r_data[34988] <= r_data[34987];
                
                r_data[34989] <= r_data[34988];
                
                r_data[34990] <= r_data[34989];
                
                r_data[34991] <= r_data[34990];
                
                r_data[34992] <= r_data[34991];
                
                r_data[34993] <= r_data[34992];
                
                r_data[34994] <= r_data[34993];
                
                r_data[34995] <= r_data[34994];
                
                r_data[34996] <= r_data[34995];
                
                r_data[34997] <= r_data[34996];
                
                r_data[34998] <= r_data[34997];
                
                r_data[34999] <= r_data[34998];
                
                r_data[35000] <= r_data[34999];
                
                r_data[35001] <= r_data[35000];
                
                r_data[35002] <= r_data[35001];
                
                r_data[35003] <= r_data[35002];
                
                r_data[35004] <= r_data[35003];
                
                r_data[35005] <= r_data[35004];
                
                r_data[35006] <= r_data[35005];
                
                r_data[35007] <= r_data[35006];
                
                r_data[35008] <= r_data[35007];
                
                r_data[35009] <= r_data[35008];
                
                r_data[35010] <= r_data[35009];
                
                r_data[35011] <= r_data[35010];
                
                r_data[35012] <= r_data[35011];
                
                r_data[35013] <= r_data[35012];
                
                r_data[35014] <= r_data[35013];
                
                r_data[35015] <= r_data[35014];
                
                r_data[35016] <= r_data[35015];
                
                r_data[35017] <= r_data[35016];
                
                r_data[35018] <= r_data[35017];
                
                r_data[35019] <= r_data[35018];
                
                r_data[35020] <= r_data[35019];
                
                r_data[35021] <= r_data[35020];
                
                r_data[35022] <= r_data[35021];
                
                r_data[35023] <= r_data[35022];
                
                r_data[35024] <= r_data[35023];
                
                r_data[35025] <= r_data[35024];
                
                r_data[35026] <= r_data[35025];
                
                r_data[35027] <= r_data[35026];
                
                r_data[35028] <= r_data[35027];
                
                r_data[35029] <= r_data[35028];
                
                r_data[35030] <= r_data[35029];
                
                r_data[35031] <= r_data[35030];
                
                r_data[35032] <= r_data[35031];
                
                r_data[35033] <= r_data[35032];
                
                r_data[35034] <= r_data[35033];
                
                r_data[35035] <= r_data[35034];
                
                r_data[35036] <= r_data[35035];
                
                r_data[35037] <= r_data[35036];
                
                r_data[35038] <= r_data[35037];
                
                r_data[35039] <= r_data[35038];
                
                r_data[35040] <= r_data[35039];
                
                r_data[35041] <= r_data[35040];
                
                r_data[35042] <= r_data[35041];
                
                r_data[35043] <= r_data[35042];
                
                r_data[35044] <= r_data[35043];
                
                r_data[35045] <= r_data[35044];
                
                r_data[35046] <= r_data[35045];
                
                r_data[35047] <= r_data[35046];
                
                r_data[35048] <= r_data[35047];
                
                r_data[35049] <= r_data[35048];
                
                r_data[35050] <= r_data[35049];
                
                r_data[35051] <= r_data[35050];
                
                r_data[35052] <= r_data[35051];
                
                r_data[35053] <= r_data[35052];
                
                r_data[35054] <= r_data[35053];
                
                r_data[35055] <= r_data[35054];
                
                r_data[35056] <= r_data[35055];
                
                r_data[35057] <= r_data[35056];
                
                r_data[35058] <= r_data[35057];
                
                r_data[35059] <= r_data[35058];
                
                r_data[35060] <= r_data[35059];
                
                r_data[35061] <= r_data[35060];
                
                r_data[35062] <= r_data[35061];
                
                r_data[35063] <= r_data[35062];
                
                r_data[35064] <= r_data[35063];
                
                r_data[35065] <= r_data[35064];
                
                r_data[35066] <= r_data[35065];
                
                r_data[35067] <= r_data[35066];
                
                r_data[35068] <= r_data[35067];
                
                r_data[35069] <= r_data[35068];
                
                r_data[35070] <= r_data[35069];
                
                r_data[35071] <= r_data[35070];
                
                r_data[35072] <= r_data[35071];
                
                r_data[35073] <= r_data[35072];
                
                r_data[35074] <= r_data[35073];
                
                r_data[35075] <= r_data[35074];
                
                r_data[35076] <= r_data[35075];
                
                r_data[35077] <= r_data[35076];
                
                r_data[35078] <= r_data[35077];
                
                r_data[35079] <= r_data[35078];
                
                r_data[35080] <= r_data[35079];
                
                r_data[35081] <= r_data[35080];
                
                r_data[35082] <= r_data[35081];
                
                r_data[35083] <= r_data[35082];
                
                r_data[35084] <= r_data[35083];
                
                r_data[35085] <= r_data[35084];
                
                r_data[35086] <= r_data[35085];
                
                r_data[35087] <= r_data[35086];
                
                r_data[35088] <= r_data[35087];
                
                r_data[35089] <= r_data[35088];
                
                r_data[35090] <= r_data[35089];
                
                r_data[35091] <= r_data[35090];
                
                r_data[35092] <= r_data[35091];
                
                r_data[35093] <= r_data[35092];
                
                r_data[35094] <= r_data[35093];
                
                r_data[35095] <= r_data[35094];
                
                r_data[35096] <= r_data[35095];
                
                r_data[35097] <= r_data[35096];
                
                r_data[35098] <= r_data[35097];
                
                r_data[35099] <= r_data[35098];
                
                r_data[35100] <= r_data[35099];
                
                r_data[35101] <= r_data[35100];
                
                r_data[35102] <= r_data[35101];
                
                r_data[35103] <= r_data[35102];
                
                r_data[35104] <= r_data[35103];
                
                r_data[35105] <= r_data[35104];
                
                r_data[35106] <= r_data[35105];
                
                r_data[35107] <= r_data[35106];
                
                r_data[35108] <= r_data[35107];
                
                r_data[35109] <= r_data[35108];
                
                r_data[35110] <= r_data[35109];
                
                r_data[35111] <= r_data[35110];
                
                r_data[35112] <= r_data[35111];
                
                r_data[35113] <= r_data[35112];
                
                r_data[35114] <= r_data[35113];
                
                r_data[35115] <= r_data[35114];
                
                r_data[35116] <= r_data[35115];
                
                r_data[35117] <= r_data[35116];
                
                r_data[35118] <= r_data[35117];
                
                r_data[35119] <= r_data[35118];
                
                r_data[35120] <= r_data[35119];
                
                r_data[35121] <= r_data[35120];
                
                r_data[35122] <= r_data[35121];
                
                r_data[35123] <= r_data[35122];
                
                r_data[35124] <= r_data[35123];
                
                r_data[35125] <= r_data[35124];
                
                r_data[35126] <= r_data[35125];
                
                r_data[35127] <= r_data[35126];
                
                r_data[35128] <= r_data[35127];
                
                r_data[35129] <= r_data[35128];
                
                r_data[35130] <= r_data[35129];
                
                r_data[35131] <= r_data[35130];
                
                r_data[35132] <= r_data[35131];
                
                r_data[35133] <= r_data[35132];
                
                r_data[35134] <= r_data[35133];
                
                r_data[35135] <= r_data[35134];
                
                r_data[35136] <= r_data[35135];
                
                r_data[35137] <= r_data[35136];
                
                r_data[35138] <= r_data[35137];
                
                r_data[35139] <= r_data[35138];
                
                r_data[35140] <= r_data[35139];
                
                r_data[35141] <= r_data[35140];
                
                r_data[35142] <= r_data[35141];
                
                r_data[35143] <= r_data[35142];
                
                r_data[35144] <= r_data[35143];
                
                r_data[35145] <= r_data[35144];
                
                r_data[35146] <= r_data[35145];
                
                r_data[35147] <= r_data[35146];
                
                r_data[35148] <= r_data[35147];
                
                r_data[35149] <= r_data[35148];
                
                r_data[35150] <= r_data[35149];
                
                r_data[35151] <= r_data[35150];
                
                r_data[35152] <= r_data[35151];
                
                r_data[35153] <= r_data[35152];
                
                r_data[35154] <= r_data[35153];
                
                r_data[35155] <= r_data[35154];
                
                r_data[35156] <= r_data[35155];
                
                r_data[35157] <= r_data[35156];
                
                r_data[35158] <= r_data[35157];
                
                r_data[35159] <= r_data[35158];
                
                r_data[35160] <= r_data[35159];
                
                r_data[35161] <= r_data[35160];
                
                r_data[35162] <= r_data[35161];
                
                r_data[35163] <= r_data[35162];
                
                r_data[35164] <= r_data[35163];
                
                r_data[35165] <= r_data[35164];
                
                r_data[35166] <= r_data[35165];
                
                r_data[35167] <= r_data[35166];
                
                r_data[35168] <= r_data[35167];
                
                r_data[35169] <= r_data[35168];
                
                r_data[35170] <= r_data[35169];
                
                r_data[35171] <= r_data[35170];
                
                r_data[35172] <= r_data[35171];
                
                r_data[35173] <= r_data[35172];
                
                r_data[35174] <= r_data[35173];
                
                r_data[35175] <= r_data[35174];
                
                r_data[35176] <= r_data[35175];
                
                r_data[35177] <= r_data[35176];
                
                r_data[35178] <= r_data[35177];
                
                r_data[35179] <= r_data[35178];
                
                r_data[35180] <= r_data[35179];
                
                r_data[35181] <= r_data[35180];
                
                r_data[35182] <= r_data[35181];
                
                r_data[35183] <= r_data[35182];
                
                r_data[35184] <= r_data[35183];
                
                r_data[35185] <= r_data[35184];
                
                r_data[35186] <= r_data[35185];
                
                r_data[35187] <= r_data[35186];
                
                r_data[35188] <= r_data[35187];
                
                r_data[35189] <= r_data[35188];
                
                r_data[35190] <= r_data[35189];
                
                r_data[35191] <= r_data[35190];
                
                r_data[35192] <= r_data[35191];
                
                r_data[35193] <= r_data[35192];
                
                r_data[35194] <= r_data[35193];
                
                r_data[35195] <= r_data[35194];
                
                r_data[35196] <= r_data[35195];
                
                r_data[35197] <= r_data[35196];
                
                r_data[35198] <= r_data[35197];
                
                r_data[35199] <= r_data[35198];
                
                r_data[35200] <= r_data[35199];
                
                r_data[35201] <= r_data[35200];
                
                r_data[35202] <= r_data[35201];
                
                r_data[35203] <= r_data[35202];
                
                r_data[35204] <= r_data[35203];
                
                r_data[35205] <= r_data[35204];
                
                r_data[35206] <= r_data[35205];
                
                r_data[35207] <= r_data[35206];
                
                r_data[35208] <= r_data[35207];
                
                r_data[35209] <= r_data[35208];
                
                r_data[35210] <= r_data[35209];
                
                r_data[35211] <= r_data[35210];
                
                r_data[35212] <= r_data[35211];
                
                r_data[35213] <= r_data[35212];
                
                r_data[35214] <= r_data[35213];
                
                r_data[35215] <= r_data[35214];
                
                r_data[35216] <= r_data[35215];
                
                r_data[35217] <= r_data[35216];
                
                r_data[35218] <= r_data[35217];
                
                r_data[35219] <= r_data[35218];
                
                r_data[35220] <= r_data[35219];
                
                r_data[35221] <= r_data[35220];
                
                r_data[35222] <= r_data[35221];
                
                r_data[35223] <= r_data[35222];
                
                r_data[35224] <= r_data[35223];
                
                r_data[35225] <= r_data[35224];
                
                r_data[35226] <= r_data[35225];
                
                r_data[35227] <= r_data[35226];
                
                r_data[35228] <= r_data[35227];
                
                r_data[35229] <= r_data[35228];
                
                r_data[35230] <= r_data[35229];
                
                r_data[35231] <= r_data[35230];
                
                r_data[35232] <= r_data[35231];
                
                r_data[35233] <= r_data[35232];
                
                r_data[35234] <= r_data[35233];
                
                r_data[35235] <= r_data[35234];
                
                r_data[35236] <= r_data[35235];
                
                r_data[35237] <= r_data[35236];
                
                r_data[35238] <= r_data[35237];
                
                r_data[35239] <= r_data[35238];
                
                r_data[35240] <= r_data[35239];
                
                r_data[35241] <= r_data[35240];
                
                r_data[35242] <= r_data[35241];
                
                r_data[35243] <= r_data[35242];
                
                r_data[35244] <= r_data[35243];
                
                r_data[35245] <= r_data[35244];
                
                r_data[35246] <= r_data[35245];
                
                r_data[35247] <= r_data[35246];
                
                r_data[35248] <= r_data[35247];
                
                r_data[35249] <= r_data[35248];
                
                r_data[35250] <= r_data[35249];
                
                r_data[35251] <= r_data[35250];
                
                r_data[35252] <= r_data[35251];
                
                r_data[35253] <= r_data[35252];
                
                r_data[35254] <= r_data[35253];
                
                r_data[35255] <= r_data[35254];
                
                r_data[35256] <= r_data[35255];
                
                r_data[35257] <= r_data[35256];
                
                r_data[35258] <= r_data[35257];
                
                r_data[35259] <= r_data[35258];
                
                r_data[35260] <= r_data[35259];
                
                r_data[35261] <= r_data[35260];
                
                r_data[35262] <= r_data[35261];
                
                r_data[35263] <= r_data[35262];
                
                r_data[35264] <= r_data[35263];
                
                r_data[35265] <= r_data[35264];
                
                r_data[35266] <= r_data[35265];
                
                r_data[35267] <= r_data[35266];
                
                r_data[35268] <= r_data[35267];
                
                r_data[35269] <= r_data[35268];
                
                r_data[35270] <= r_data[35269];
                
                r_data[35271] <= r_data[35270];
                
                r_data[35272] <= r_data[35271];
                
                r_data[35273] <= r_data[35272];
                
                r_data[35274] <= r_data[35273];
                
                r_data[35275] <= r_data[35274];
                
                r_data[35276] <= r_data[35275];
                
                r_data[35277] <= r_data[35276];
                
                r_data[35278] <= r_data[35277];
                
                r_data[35279] <= r_data[35278];
                
                r_data[35280] <= r_data[35279];
                
                r_data[35281] <= r_data[35280];
                
                r_data[35282] <= r_data[35281];
                
                r_data[35283] <= r_data[35282];
                
                r_data[35284] <= r_data[35283];
                
                r_data[35285] <= r_data[35284];
                
                r_data[35286] <= r_data[35285];
                
                r_data[35287] <= r_data[35286];
                
                r_data[35288] <= r_data[35287];
                
                r_data[35289] <= r_data[35288];
                
                r_data[35290] <= r_data[35289];
                
                r_data[35291] <= r_data[35290];
                
                r_data[35292] <= r_data[35291];
                
                r_data[35293] <= r_data[35292];
                
                r_data[35294] <= r_data[35293];
                
                r_data[35295] <= r_data[35294];
                
                r_data[35296] <= r_data[35295];
                
                r_data[35297] <= r_data[35296];
                
                r_data[35298] <= r_data[35297];
                
                r_data[35299] <= r_data[35298];
                
                r_data[35300] <= r_data[35299];
                
                r_data[35301] <= r_data[35300];
                
                r_data[35302] <= r_data[35301];
                
                r_data[35303] <= r_data[35302];
                
                r_data[35304] <= r_data[35303];
                
                r_data[35305] <= r_data[35304];
                
                r_data[35306] <= r_data[35305];
                
                r_data[35307] <= r_data[35306];
                
                r_data[35308] <= r_data[35307];
                
                r_data[35309] <= r_data[35308];
                
                r_data[35310] <= r_data[35309];
                
                r_data[35311] <= r_data[35310];
                
                r_data[35312] <= r_data[35311];
                
                r_data[35313] <= r_data[35312];
                
                r_data[35314] <= r_data[35313];
                
                r_data[35315] <= r_data[35314];
                
                r_data[35316] <= r_data[35315];
                
                r_data[35317] <= r_data[35316];
                
                r_data[35318] <= r_data[35317];
                
                r_data[35319] <= r_data[35318];
                
                r_data[35320] <= r_data[35319];
                
                r_data[35321] <= r_data[35320];
                
                r_data[35322] <= r_data[35321];
                
                r_data[35323] <= r_data[35322];
                
                r_data[35324] <= r_data[35323];
                
                r_data[35325] <= r_data[35324];
                
                r_data[35326] <= r_data[35325];
                
                r_data[35327] <= r_data[35326];
                
                r_data[35328] <= r_data[35327];
                
                r_data[35329] <= r_data[35328];
                
                r_data[35330] <= r_data[35329];
                
                r_data[35331] <= r_data[35330];
                
                r_data[35332] <= r_data[35331];
                
                r_data[35333] <= r_data[35332];
                
                r_data[35334] <= r_data[35333];
                
                r_data[35335] <= r_data[35334];
                
                r_data[35336] <= r_data[35335];
                
                r_data[35337] <= r_data[35336];
                
                r_data[35338] <= r_data[35337];
                
                r_data[35339] <= r_data[35338];
                
                r_data[35340] <= r_data[35339];
                
                r_data[35341] <= r_data[35340];
                
                r_data[35342] <= r_data[35341];
                
                r_data[35343] <= r_data[35342];
                
                r_data[35344] <= r_data[35343];
                
                r_data[35345] <= r_data[35344];
                
                r_data[35346] <= r_data[35345];
                
                r_data[35347] <= r_data[35346];
                
                r_data[35348] <= r_data[35347];
                
                r_data[35349] <= r_data[35348];
                
                r_data[35350] <= r_data[35349];
                
                r_data[35351] <= r_data[35350];
                
                r_data[35352] <= r_data[35351];
                
                r_data[35353] <= r_data[35352];
                
                r_data[35354] <= r_data[35353];
                
                r_data[35355] <= r_data[35354];
                
                r_data[35356] <= r_data[35355];
                
                r_data[35357] <= r_data[35356];
                
                r_data[35358] <= r_data[35357];
                
                r_data[35359] <= r_data[35358];
                
                r_data[35360] <= r_data[35359];
                
                r_data[35361] <= r_data[35360];
                
                r_data[35362] <= r_data[35361];
                
                r_data[35363] <= r_data[35362];
                
                r_data[35364] <= r_data[35363];
                
                r_data[35365] <= r_data[35364];
                
                r_data[35366] <= r_data[35365];
                
                r_data[35367] <= r_data[35366];
                
                r_data[35368] <= r_data[35367];
                
                r_data[35369] <= r_data[35368];
                
                r_data[35370] <= r_data[35369];
                
                r_data[35371] <= r_data[35370];
                
                r_data[35372] <= r_data[35371];
                
                r_data[35373] <= r_data[35372];
                
                r_data[35374] <= r_data[35373];
                
                r_data[35375] <= r_data[35374];
                
                r_data[35376] <= r_data[35375];
                
                r_data[35377] <= r_data[35376];
                
                r_data[35378] <= r_data[35377];
                
                r_data[35379] <= r_data[35378];
                
                r_data[35380] <= r_data[35379];
                
                r_data[35381] <= r_data[35380];
                
                r_data[35382] <= r_data[35381];
                
                r_data[35383] <= r_data[35382];
                
                r_data[35384] <= r_data[35383];
                
                r_data[35385] <= r_data[35384];
                
                r_data[35386] <= r_data[35385];
                
                r_data[35387] <= r_data[35386];
                
                r_data[35388] <= r_data[35387];
                
                r_data[35389] <= r_data[35388];
                
                r_data[35390] <= r_data[35389];
                
                r_data[35391] <= r_data[35390];
                
                r_data[35392] <= r_data[35391];
                
                r_data[35393] <= r_data[35392];
                
                r_data[35394] <= r_data[35393];
                
                r_data[35395] <= r_data[35394];
                
                r_data[35396] <= r_data[35395];
                
                r_data[35397] <= r_data[35396];
                
                r_data[35398] <= r_data[35397];
                
                r_data[35399] <= r_data[35398];
                
                r_data[35400] <= r_data[35399];
                
                r_data[35401] <= r_data[35400];
                
                r_data[35402] <= r_data[35401];
                
                r_data[35403] <= r_data[35402];
                
                r_data[35404] <= r_data[35403];
                
                r_data[35405] <= r_data[35404];
                
                r_data[35406] <= r_data[35405];
                
                r_data[35407] <= r_data[35406];
                
                r_data[35408] <= r_data[35407];
                
                r_data[35409] <= r_data[35408];
                
                r_data[35410] <= r_data[35409];
                
                r_data[35411] <= r_data[35410];
                
                r_data[35412] <= r_data[35411];
                
                r_data[35413] <= r_data[35412];
                
                r_data[35414] <= r_data[35413];
                
                r_data[35415] <= r_data[35414];
                
                r_data[35416] <= r_data[35415];
                
                r_data[35417] <= r_data[35416];
                
                r_data[35418] <= r_data[35417];
                
                r_data[35419] <= r_data[35418];
                
                r_data[35420] <= r_data[35419];
                
                r_data[35421] <= r_data[35420];
                
                r_data[35422] <= r_data[35421];
                
                r_data[35423] <= r_data[35422];
                
                r_data[35424] <= r_data[35423];
                
                r_data[35425] <= r_data[35424];
                
                r_data[35426] <= r_data[35425];
                
                r_data[35427] <= r_data[35426];
                
                r_data[35428] <= r_data[35427];
                
                r_data[35429] <= r_data[35428];
                
                r_data[35430] <= r_data[35429];
                
                r_data[35431] <= r_data[35430];
                
                r_data[35432] <= r_data[35431];
                
                r_data[35433] <= r_data[35432];
                
                r_data[35434] <= r_data[35433];
                
                r_data[35435] <= r_data[35434];
                
                r_data[35436] <= r_data[35435];
                
                r_data[35437] <= r_data[35436];
                
                r_data[35438] <= r_data[35437];
                
                r_data[35439] <= r_data[35438];
                
                r_data[35440] <= r_data[35439];
                
                r_data[35441] <= r_data[35440];
                
                r_data[35442] <= r_data[35441];
                
                r_data[35443] <= r_data[35442];
                
                r_data[35444] <= r_data[35443];
                
                r_data[35445] <= r_data[35444];
                
                r_data[35446] <= r_data[35445];
                
                r_data[35447] <= r_data[35446];
                
                r_data[35448] <= r_data[35447];
                
                r_data[35449] <= r_data[35448];
                
                r_data[35450] <= r_data[35449];
                
                r_data[35451] <= r_data[35450];
                
                r_data[35452] <= r_data[35451];
                
                r_data[35453] <= r_data[35452];
                
                r_data[35454] <= r_data[35453];
                
                r_data[35455] <= r_data[35454];
                
                r_data[35456] <= r_data[35455];
                
                r_data[35457] <= r_data[35456];
                
                r_data[35458] <= r_data[35457];
                
                r_data[35459] <= r_data[35458];
                
                r_data[35460] <= r_data[35459];
                
                r_data[35461] <= r_data[35460];
                
                r_data[35462] <= r_data[35461];
                
                r_data[35463] <= r_data[35462];
                
                r_data[35464] <= r_data[35463];
                
                r_data[35465] <= r_data[35464];
                
                r_data[35466] <= r_data[35465];
                
                r_data[35467] <= r_data[35466];
                
                r_data[35468] <= r_data[35467];
                
                r_data[35469] <= r_data[35468];
                
                r_data[35470] <= r_data[35469];
                
                r_data[35471] <= r_data[35470];
                
                r_data[35472] <= r_data[35471];
                
                r_data[35473] <= r_data[35472];
                
                r_data[35474] <= r_data[35473];
                
                r_data[35475] <= r_data[35474];
                
                r_data[35476] <= r_data[35475];
                
                r_data[35477] <= r_data[35476];
                
                r_data[35478] <= r_data[35477];
                
                r_data[35479] <= r_data[35478];
                
                r_data[35480] <= r_data[35479];
                
                r_data[35481] <= r_data[35480];
                
                r_data[35482] <= r_data[35481];
                
                r_data[35483] <= r_data[35482];
                
                r_data[35484] <= r_data[35483];
                
                r_data[35485] <= r_data[35484];
                
                r_data[35486] <= r_data[35485];
                
                r_data[35487] <= r_data[35486];
                
                r_data[35488] <= r_data[35487];
                
                r_data[35489] <= r_data[35488];
                
                r_data[35490] <= r_data[35489];
                
                r_data[35491] <= r_data[35490];
                
                r_data[35492] <= r_data[35491];
                
                r_data[35493] <= r_data[35492];
                
                r_data[35494] <= r_data[35493];
                
                r_data[35495] <= r_data[35494];
                
                r_data[35496] <= r_data[35495];
                
                r_data[35497] <= r_data[35496];
                
                r_data[35498] <= r_data[35497];
                
                r_data[35499] <= r_data[35498];
                
                r_data[35500] <= r_data[35499];
                
                r_data[35501] <= r_data[35500];
                
                r_data[35502] <= r_data[35501];
                
                r_data[35503] <= r_data[35502];
                
                r_data[35504] <= r_data[35503];
                
                r_data[35505] <= r_data[35504];
                
                r_data[35506] <= r_data[35505];
                
                r_data[35507] <= r_data[35506];
                
                r_data[35508] <= r_data[35507];
                
                r_data[35509] <= r_data[35508];
                
                r_data[35510] <= r_data[35509];
                
                r_data[35511] <= r_data[35510];
                
                r_data[35512] <= r_data[35511];
                
                r_data[35513] <= r_data[35512];
                
                r_data[35514] <= r_data[35513];
                
                r_data[35515] <= r_data[35514];
                
                r_data[35516] <= r_data[35515];
                
                r_data[35517] <= r_data[35516];
                
                r_data[35518] <= r_data[35517];
                
                r_data[35519] <= r_data[35518];
                
                r_data[35520] <= r_data[35519];
                
                r_data[35521] <= r_data[35520];
                
                r_data[35522] <= r_data[35521];
                
                r_data[35523] <= r_data[35522];
                
                r_data[35524] <= r_data[35523];
                
                r_data[35525] <= r_data[35524];
                
                r_data[35526] <= r_data[35525];
                
                r_data[35527] <= r_data[35526];
                
                r_data[35528] <= r_data[35527];
                
                r_data[35529] <= r_data[35528];
                
                r_data[35530] <= r_data[35529];
                
                r_data[35531] <= r_data[35530];
                
                r_data[35532] <= r_data[35531];
                
                r_data[35533] <= r_data[35532];
                
                r_data[35534] <= r_data[35533];
                
                r_data[35535] <= r_data[35534];
                
                r_data[35536] <= r_data[35535];
                
                r_data[35537] <= r_data[35536];
                
                r_data[35538] <= r_data[35537];
                
                r_data[35539] <= r_data[35538];
                
                r_data[35540] <= r_data[35539];
                
                r_data[35541] <= r_data[35540];
                
                r_data[35542] <= r_data[35541];
                
                r_data[35543] <= r_data[35542];
                
                r_data[35544] <= r_data[35543];
                
                r_data[35545] <= r_data[35544];
                
                r_data[35546] <= r_data[35545];
                
                r_data[35547] <= r_data[35546];
                
                r_data[35548] <= r_data[35547];
                
                r_data[35549] <= r_data[35548];
                
                r_data[35550] <= r_data[35549];
                
                r_data[35551] <= r_data[35550];
                
                r_data[35552] <= r_data[35551];
                
                r_data[35553] <= r_data[35552];
                
                r_data[35554] <= r_data[35553];
                
                r_data[35555] <= r_data[35554];
                
                r_data[35556] <= r_data[35555];
                
                r_data[35557] <= r_data[35556];
                
                r_data[35558] <= r_data[35557];
                
                r_data[35559] <= r_data[35558];
                
                r_data[35560] <= r_data[35559];
                
                r_data[35561] <= r_data[35560];
                
                r_data[35562] <= r_data[35561];
                
                r_data[35563] <= r_data[35562];
                
                r_data[35564] <= r_data[35563];
                
                r_data[35565] <= r_data[35564];
                
                r_data[35566] <= r_data[35565];
                
                r_data[35567] <= r_data[35566];
                
                r_data[35568] <= r_data[35567];
                
                r_data[35569] <= r_data[35568];
                
                r_data[35570] <= r_data[35569];
                
                r_data[35571] <= r_data[35570];
                
                r_data[35572] <= r_data[35571];
                
                r_data[35573] <= r_data[35572];
                
                r_data[35574] <= r_data[35573];
                
                r_data[35575] <= r_data[35574];
                
                r_data[35576] <= r_data[35575];
                
                r_data[35577] <= r_data[35576];
                
                r_data[35578] <= r_data[35577];
                
                r_data[35579] <= r_data[35578];
                
                r_data[35580] <= r_data[35579];
                
                r_data[35581] <= r_data[35580];
                
                r_data[35582] <= r_data[35581];
                
                r_data[35583] <= r_data[35582];
                
                r_data[35584] <= r_data[35583];
                
                r_data[35585] <= r_data[35584];
                
                r_data[35586] <= r_data[35585];
                
                r_data[35587] <= r_data[35586];
                
                r_data[35588] <= r_data[35587];
                
                r_data[35589] <= r_data[35588];
                
                r_data[35590] <= r_data[35589];
                
                r_data[35591] <= r_data[35590];
                
                r_data[35592] <= r_data[35591];
                
                r_data[35593] <= r_data[35592];
                
                r_data[35594] <= r_data[35593];
                
                r_data[35595] <= r_data[35594];
                
                r_data[35596] <= r_data[35595];
                
                r_data[35597] <= r_data[35596];
                
                r_data[35598] <= r_data[35597];
                
                r_data[35599] <= r_data[35598];
                
                r_data[35600] <= r_data[35599];
                
                r_data[35601] <= r_data[35600];
                
                r_data[35602] <= r_data[35601];
                
                r_data[35603] <= r_data[35602];
                
                r_data[35604] <= r_data[35603];
                
                r_data[35605] <= r_data[35604];
                
                r_data[35606] <= r_data[35605];
                
                r_data[35607] <= r_data[35606];
                
                r_data[35608] <= r_data[35607];
                
                r_data[35609] <= r_data[35608];
                
                r_data[35610] <= r_data[35609];
                
                r_data[35611] <= r_data[35610];
                
                r_data[35612] <= r_data[35611];
                
                r_data[35613] <= r_data[35612];
                
                r_data[35614] <= r_data[35613];
                
                r_data[35615] <= r_data[35614];
                
                r_data[35616] <= r_data[35615];
                
                r_data[35617] <= r_data[35616];
                
                r_data[35618] <= r_data[35617];
                
                r_data[35619] <= r_data[35618];
                
                r_data[35620] <= r_data[35619];
                
                r_data[35621] <= r_data[35620];
                
                r_data[35622] <= r_data[35621];
                
                r_data[35623] <= r_data[35622];
                
                r_data[35624] <= r_data[35623];
                
                r_data[35625] <= r_data[35624];
                
                r_data[35626] <= r_data[35625];
                
                r_data[35627] <= r_data[35626];
                
                r_data[35628] <= r_data[35627];
                
                r_data[35629] <= r_data[35628];
                
                r_data[35630] <= r_data[35629];
                
                r_data[35631] <= r_data[35630];
                
                r_data[35632] <= r_data[35631];
                
                r_data[35633] <= r_data[35632];
                
                r_data[35634] <= r_data[35633];
                
                r_data[35635] <= r_data[35634];
                
                r_data[35636] <= r_data[35635];
                
                r_data[35637] <= r_data[35636];
                
                r_data[35638] <= r_data[35637];
                
                r_data[35639] <= r_data[35638];
                
                r_data[35640] <= r_data[35639];
                
                r_data[35641] <= r_data[35640];
                
                r_data[35642] <= r_data[35641];
                
                r_data[35643] <= r_data[35642];
                
                r_data[35644] <= r_data[35643];
                
                r_data[35645] <= r_data[35644];
                
                r_data[35646] <= r_data[35645];
                
                r_data[35647] <= r_data[35646];
                
                r_data[35648] <= r_data[35647];
                
                r_data[35649] <= r_data[35648];
                
                r_data[35650] <= r_data[35649];
                
                r_data[35651] <= r_data[35650];
                
                r_data[35652] <= r_data[35651];
                
                r_data[35653] <= r_data[35652];
                
                r_data[35654] <= r_data[35653];
                
                r_data[35655] <= r_data[35654];
                
                r_data[35656] <= r_data[35655];
                
                r_data[35657] <= r_data[35656];
                
                r_data[35658] <= r_data[35657];
                
                r_data[35659] <= r_data[35658];
                
                r_data[35660] <= r_data[35659];
                
                r_data[35661] <= r_data[35660];
                
                r_data[35662] <= r_data[35661];
                
                r_data[35663] <= r_data[35662];
                
                r_data[35664] <= r_data[35663];
                
                r_data[35665] <= r_data[35664];
                
                r_data[35666] <= r_data[35665];
                
                r_data[35667] <= r_data[35666];
                
                r_data[35668] <= r_data[35667];
                
                r_data[35669] <= r_data[35668];
                
                r_data[35670] <= r_data[35669];
                
                r_data[35671] <= r_data[35670];
                
                r_data[35672] <= r_data[35671];
                
                r_data[35673] <= r_data[35672];
                
                r_data[35674] <= r_data[35673];
                
                r_data[35675] <= r_data[35674];
                
                r_data[35676] <= r_data[35675];
                
                r_data[35677] <= r_data[35676];
                
                r_data[35678] <= r_data[35677];
                
                r_data[35679] <= r_data[35678];
                
                r_data[35680] <= r_data[35679];
                
                r_data[35681] <= r_data[35680];
                
                r_data[35682] <= r_data[35681];
                
                r_data[35683] <= r_data[35682];
                
                r_data[35684] <= r_data[35683];
                
                r_data[35685] <= r_data[35684];
                
                r_data[35686] <= r_data[35685];
                
                r_data[35687] <= r_data[35686];
                
                r_data[35688] <= r_data[35687];
                
                r_data[35689] <= r_data[35688];
                
                r_data[35690] <= r_data[35689];
                
                r_data[35691] <= r_data[35690];
                
                r_data[35692] <= r_data[35691];
                
                r_data[35693] <= r_data[35692];
                
                r_data[35694] <= r_data[35693];
                
                r_data[35695] <= r_data[35694];
                
                r_data[35696] <= r_data[35695];
                
                r_data[35697] <= r_data[35696];
                
                r_data[35698] <= r_data[35697];
                
                r_data[35699] <= r_data[35698];
                
                r_data[35700] <= r_data[35699];
                
                r_data[35701] <= r_data[35700];
                
                r_data[35702] <= r_data[35701];
                
                r_data[35703] <= r_data[35702];
                
                r_data[35704] <= r_data[35703];
                
                r_data[35705] <= r_data[35704];
                
                r_data[35706] <= r_data[35705];
                
                r_data[35707] <= r_data[35706];
                
                r_data[35708] <= r_data[35707];
                
                r_data[35709] <= r_data[35708];
                
                r_data[35710] <= r_data[35709];
                
                r_data[35711] <= r_data[35710];
                
                r_data[35712] <= r_data[35711];
                
                r_data[35713] <= r_data[35712];
                
                r_data[35714] <= r_data[35713];
                
                r_data[35715] <= r_data[35714];
                
                r_data[35716] <= r_data[35715];
                
                r_data[35717] <= r_data[35716];
                
                r_data[35718] <= r_data[35717];
                
                r_data[35719] <= r_data[35718];
                
                r_data[35720] <= r_data[35719];
                
                r_data[35721] <= r_data[35720];
                
                r_data[35722] <= r_data[35721];
                
                r_data[35723] <= r_data[35722];
                
                r_data[35724] <= r_data[35723];
                
                r_data[35725] <= r_data[35724];
                
                r_data[35726] <= r_data[35725];
                
                r_data[35727] <= r_data[35726];
                
                r_data[35728] <= r_data[35727];
                
                r_data[35729] <= r_data[35728];
                
                r_data[35730] <= r_data[35729];
                
                r_data[35731] <= r_data[35730];
                
                r_data[35732] <= r_data[35731];
                
                r_data[35733] <= r_data[35732];
                
                r_data[35734] <= r_data[35733];
                
                r_data[35735] <= r_data[35734];
                
                r_data[35736] <= r_data[35735];
                
                r_data[35737] <= r_data[35736];
                
                r_data[35738] <= r_data[35737];
                
                r_data[35739] <= r_data[35738];
                
                r_data[35740] <= r_data[35739];
                
                r_data[35741] <= r_data[35740];
                
                r_data[35742] <= r_data[35741];
                
                r_data[35743] <= r_data[35742];
                
                r_data[35744] <= r_data[35743];
                
                r_data[35745] <= r_data[35744];
                
                r_data[35746] <= r_data[35745];
                
                r_data[35747] <= r_data[35746];
                
                r_data[35748] <= r_data[35747];
                
                r_data[35749] <= r_data[35748];
                
                r_data[35750] <= r_data[35749];
                
                r_data[35751] <= r_data[35750];
                
                r_data[35752] <= r_data[35751];
                
                r_data[35753] <= r_data[35752];
                
                r_data[35754] <= r_data[35753];
                
                r_data[35755] <= r_data[35754];
                
                r_data[35756] <= r_data[35755];
                
                r_data[35757] <= r_data[35756];
                
                r_data[35758] <= r_data[35757];
                
                r_data[35759] <= r_data[35758];
                
                r_data[35760] <= r_data[35759];
                
                r_data[35761] <= r_data[35760];
                
                r_data[35762] <= r_data[35761];
                
                r_data[35763] <= r_data[35762];
                
                r_data[35764] <= r_data[35763];
                
                r_data[35765] <= r_data[35764];
                
                r_data[35766] <= r_data[35765];
                
                r_data[35767] <= r_data[35766];
                
                r_data[35768] <= r_data[35767];
                
                r_data[35769] <= r_data[35768];
                
                r_data[35770] <= r_data[35769];
                
                r_data[35771] <= r_data[35770];
                
                r_data[35772] <= r_data[35771];
                
                r_data[35773] <= r_data[35772];
                
                r_data[35774] <= r_data[35773];
                
                r_data[35775] <= r_data[35774];
                
                r_data[35776] <= r_data[35775];
                
                r_data[35777] <= r_data[35776];
                
                r_data[35778] <= r_data[35777];
                
                r_data[35779] <= r_data[35778];
                
                r_data[35780] <= r_data[35779];
                
                r_data[35781] <= r_data[35780];
                
                r_data[35782] <= r_data[35781];
                
                r_data[35783] <= r_data[35782];
                
                r_data[35784] <= r_data[35783];
                
                r_data[35785] <= r_data[35784];
                
                r_data[35786] <= r_data[35785];
                
                r_data[35787] <= r_data[35786];
                
                r_data[35788] <= r_data[35787];
                
                r_data[35789] <= r_data[35788];
                
                r_data[35790] <= r_data[35789];
                
                r_data[35791] <= r_data[35790];
                
                r_data[35792] <= r_data[35791];
                
                r_data[35793] <= r_data[35792];
                
                r_data[35794] <= r_data[35793];
                
                r_data[35795] <= r_data[35794];
                
                r_data[35796] <= r_data[35795];
                
                r_data[35797] <= r_data[35796];
                
                r_data[35798] <= r_data[35797];
                
                r_data[35799] <= r_data[35798];
                
                r_data[35800] <= r_data[35799];
                
                r_data[35801] <= r_data[35800];
                
                r_data[35802] <= r_data[35801];
                
                r_data[35803] <= r_data[35802];
                
                r_data[35804] <= r_data[35803];
                
                r_data[35805] <= r_data[35804];
                
                r_data[35806] <= r_data[35805];
                
                r_data[35807] <= r_data[35806];
                
                r_data[35808] <= r_data[35807];
                
                r_data[35809] <= r_data[35808];
                
                r_data[35810] <= r_data[35809];
                
                r_data[35811] <= r_data[35810];
                
                r_data[35812] <= r_data[35811];
                
                r_data[35813] <= r_data[35812];
                
                r_data[35814] <= r_data[35813];
                
                r_data[35815] <= r_data[35814];
                
                r_data[35816] <= r_data[35815];
                
                r_data[35817] <= r_data[35816];
                
                r_data[35818] <= r_data[35817];
                
                r_data[35819] <= r_data[35818];
                
                r_data[35820] <= r_data[35819];
                
                r_data[35821] <= r_data[35820];
                
                r_data[35822] <= r_data[35821];
                
                r_data[35823] <= r_data[35822];
                
                r_data[35824] <= r_data[35823];
                
                r_data[35825] <= r_data[35824];
                
                r_data[35826] <= r_data[35825];
                
                r_data[35827] <= r_data[35826];
                
                r_data[35828] <= r_data[35827];
                
                r_data[35829] <= r_data[35828];
                
                r_data[35830] <= r_data[35829];
                
                r_data[35831] <= r_data[35830];
                
                r_data[35832] <= r_data[35831];
                
                r_data[35833] <= r_data[35832];
                
                r_data[35834] <= r_data[35833];
                
                r_data[35835] <= r_data[35834];
                
                r_data[35836] <= r_data[35835];
                
                r_data[35837] <= r_data[35836];
                
                r_data[35838] <= r_data[35837];
                
                r_data[35839] <= r_data[35838];
                
                r_data[35840] <= r_data[35839];
                
                r_data[35841] <= r_data[35840];
                
                r_data[35842] <= r_data[35841];
                
                r_data[35843] <= r_data[35842];
                
                r_data[35844] <= r_data[35843];
                
                r_data[35845] <= r_data[35844];
                
                r_data[35846] <= r_data[35845];
                
                r_data[35847] <= r_data[35846];
                
                r_data[35848] <= r_data[35847];
                
                r_data[35849] <= r_data[35848];
                
                r_data[35850] <= r_data[35849];
                
                r_data[35851] <= r_data[35850];
                
                r_data[35852] <= r_data[35851];
                
                r_data[35853] <= r_data[35852];
                
                r_data[35854] <= r_data[35853];
                
                r_data[35855] <= r_data[35854];
                
                r_data[35856] <= r_data[35855];
                
                r_data[35857] <= r_data[35856];
                
                r_data[35858] <= r_data[35857];
                
                r_data[35859] <= r_data[35858];
                
                r_data[35860] <= r_data[35859];
                
                r_data[35861] <= r_data[35860];
                
                r_data[35862] <= r_data[35861];
                
                r_data[35863] <= r_data[35862];
                
                r_data[35864] <= r_data[35863];
                
                r_data[35865] <= r_data[35864];
                
                r_data[35866] <= r_data[35865];
                
                r_data[35867] <= r_data[35866];
                
                r_data[35868] <= r_data[35867];
                
                r_data[35869] <= r_data[35868];
                
                r_data[35870] <= r_data[35869];
                
                r_data[35871] <= r_data[35870];
                
                r_data[35872] <= r_data[35871];
                
                r_data[35873] <= r_data[35872];
                
                r_data[35874] <= r_data[35873];
                
                r_data[35875] <= r_data[35874];
                
                r_data[35876] <= r_data[35875];
                
                r_data[35877] <= r_data[35876];
                
                r_data[35878] <= r_data[35877];
                
                r_data[35879] <= r_data[35878];
                
                r_data[35880] <= r_data[35879];
                
                r_data[35881] <= r_data[35880];
                
                r_data[35882] <= r_data[35881];
                
                r_data[35883] <= r_data[35882];
                
                r_data[35884] <= r_data[35883];
                
                r_data[35885] <= r_data[35884];
                
                r_data[35886] <= r_data[35885];
                
                r_data[35887] <= r_data[35886];
                
                r_data[35888] <= r_data[35887];
                
                r_data[35889] <= r_data[35888];
                
                r_data[35890] <= r_data[35889];
                
                r_data[35891] <= r_data[35890];
                
                r_data[35892] <= r_data[35891];
                
                r_data[35893] <= r_data[35892];
                
                r_data[35894] <= r_data[35893];
                
                r_data[35895] <= r_data[35894];
                
                r_data[35896] <= r_data[35895];
                
                r_data[35897] <= r_data[35896];
                
                r_data[35898] <= r_data[35897];
                
                r_data[35899] <= r_data[35898];
                
                r_data[35900] <= r_data[35899];
                
                r_data[35901] <= r_data[35900];
                
                r_data[35902] <= r_data[35901];
                
                r_data[35903] <= r_data[35902];
                
                r_data[35904] <= r_data[35903];
                
                r_data[35905] <= r_data[35904];
                
                r_data[35906] <= r_data[35905];
                
                r_data[35907] <= r_data[35906];
                
                r_data[35908] <= r_data[35907];
                
                r_data[35909] <= r_data[35908];
                
                r_data[35910] <= r_data[35909];
                
                r_data[35911] <= r_data[35910];
                
                r_data[35912] <= r_data[35911];
                
                r_data[35913] <= r_data[35912];
                
                r_data[35914] <= r_data[35913];
                
                r_data[35915] <= r_data[35914];
                
                r_data[35916] <= r_data[35915];
                
                r_data[35917] <= r_data[35916];
                
                r_data[35918] <= r_data[35917];
                
                r_data[35919] <= r_data[35918];
                
                r_data[35920] <= r_data[35919];
                
                r_data[35921] <= r_data[35920];
                
                r_data[35922] <= r_data[35921];
                
                r_data[35923] <= r_data[35922];
                
                r_data[35924] <= r_data[35923];
                
                r_data[35925] <= r_data[35924];
                
                r_data[35926] <= r_data[35925];
                
                r_data[35927] <= r_data[35926];
                
                r_data[35928] <= r_data[35927];
                
                r_data[35929] <= r_data[35928];
                
                r_data[35930] <= r_data[35929];
                
                r_data[35931] <= r_data[35930];
                
                r_data[35932] <= r_data[35931];
                
                r_data[35933] <= r_data[35932];
                
                r_data[35934] <= r_data[35933];
                
                r_data[35935] <= r_data[35934];
                
                r_data[35936] <= r_data[35935];
                
                r_data[35937] <= r_data[35936];
                
                r_data[35938] <= r_data[35937];
                
                r_data[35939] <= r_data[35938];
                
                r_data[35940] <= r_data[35939];
                
                r_data[35941] <= r_data[35940];
                
                r_data[35942] <= r_data[35941];
                
                r_data[35943] <= r_data[35942];
                
                r_data[35944] <= r_data[35943];
                
                r_data[35945] <= r_data[35944];
                
                r_data[35946] <= r_data[35945];
                
                r_data[35947] <= r_data[35946];
                
                r_data[35948] <= r_data[35947];
                
                r_data[35949] <= r_data[35948];
                
                r_data[35950] <= r_data[35949];
                
                r_data[35951] <= r_data[35950];
                
                r_data[35952] <= r_data[35951];
                
                r_data[35953] <= r_data[35952];
                
                r_data[35954] <= r_data[35953];
                
                r_data[35955] <= r_data[35954];
                
                r_data[35956] <= r_data[35955];
                
                r_data[35957] <= r_data[35956];
                
                r_data[35958] <= r_data[35957];
                
                r_data[35959] <= r_data[35958];
                
                r_data[35960] <= r_data[35959];
                
                r_data[35961] <= r_data[35960];
                
                r_data[35962] <= r_data[35961];
                
                r_data[35963] <= r_data[35962];
                
                r_data[35964] <= r_data[35963];
                
                r_data[35965] <= r_data[35964];
                
                r_data[35966] <= r_data[35965];
                
                r_data[35967] <= r_data[35966];
                
                r_data[35968] <= r_data[35967];
                
                r_data[35969] <= r_data[35968];
                
                r_data[35970] <= r_data[35969];
                
                r_data[35971] <= r_data[35970];
                
                r_data[35972] <= r_data[35971];
                
                r_data[35973] <= r_data[35972];
                
                r_data[35974] <= r_data[35973];
                
                r_data[35975] <= r_data[35974];
                
                r_data[35976] <= r_data[35975];
                
                r_data[35977] <= r_data[35976];
                
                r_data[35978] <= r_data[35977];
                
                r_data[35979] <= r_data[35978];
                
                r_data[35980] <= r_data[35979];
                
                r_data[35981] <= r_data[35980];
                
                r_data[35982] <= r_data[35981];
                
                r_data[35983] <= r_data[35982];
                
                r_data[35984] <= r_data[35983];
                
                r_data[35985] <= r_data[35984];
                
                r_data[35986] <= r_data[35985];
                
                r_data[35987] <= r_data[35986];
                
                r_data[35988] <= r_data[35987];
                
                r_data[35989] <= r_data[35988];
                
                r_data[35990] <= r_data[35989];
                
                r_data[35991] <= r_data[35990];
                
                r_data[35992] <= r_data[35991];
                
                r_data[35993] <= r_data[35992];
                
                r_data[35994] <= r_data[35993];
                
                r_data[35995] <= r_data[35994];
                
                r_data[35996] <= r_data[35995];
                
                r_data[35997] <= r_data[35996];
                
                r_data[35998] <= r_data[35997];
                
                r_data[35999] <= r_data[35998];
                
                r_data[36000] <= r_data[35999];
                
                r_data[36001] <= r_data[36000];
                
                r_data[36002] <= r_data[36001];
                
                r_data[36003] <= r_data[36002];
                
                r_data[36004] <= r_data[36003];
                
                r_data[36005] <= r_data[36004];
                
                r_data[36006] <= r_data[36005];
                
                r_data[36007] <= r_data[36006];
                
                r_data[36008] <= r_data[36007];
                
                r_data[36009] <= r_data[36008];
                
                r_data[36010] <= r_data[36009];
                
                r_data[36011] <= r_data[36010];
                
                r_data[36012] <= r_data[36011];
                
                r_data[36013] <= r_data[36012];
                
                r_data[36014] <= r_data[36013];
                
                r_data[36015] <= r_data[36014];
                
                r_data[36016] <= r_data[36015];
                
                r_data[36017] <= r_data[36016];
                
                r_data[36018] <= r_data[36017];
                
                r_data[36019] <= r_data[36018];
                
                r_data[36020] <= r_data[36019];
                
                r_data[36021] <= r_data[36020];
                
                r_data[36022] <= r_data[36021];
                
                r_data[36023] <= r_data[36022];
                
                r_data[36024] <= r_data[36023];
                
                r_data[36025] <= r_data[36024];
                
                r_data[36026] <= r_data[36025];
                
                r_data[36027] <= r_data[36026];
                
                r_data[36028] <= r_data[36027];
                
                r_data[36029] <= r_data[36028];
                
                r_data[36030] <= r_data[36029];
                
                r_data[36031] <= r_data[36030];
                
                r_data[36032] <= r_data[36031];
                
                r_data[36033] <= r_data[36032];
                
                r_data[36034] <= r_data[36033];
                
                r_data[36035] <= r_data[36034];
                
                r_data[36036] <= r_data[36035];
                
                r_data[36037] <= r_data[36036];
                
                r_data[36038] <= r_data[36037];
                
                r_data[36039] <= r_data[36038];
                
                r_data[36040] <= r_data[36039];
                
                r_data[36041] <= r_data[36040];
                
                r_data[36042] <= r_data[36041];
                
                r_data[36043] <= r_data[36042];
                
                r_data[36044] <= r_data[36043];
                
                r_data[36045] <= r_data[36044];
                
                r_data[36046] <= r_data[36045];
                
                r_data[36047] <= r_data[36046];
                
                r_data[36048] <= r_data[36047];
                
                r_data[36049] <= r_data[36048];
                
                r_data[36050] <= r_data[36049];
                
                r_data[36051] <= r_data[36050];
                
                r_data[36052] <= r_data[36051];
                
                r_data[36053] <= r_data[36052];
                
                r_data[36054] <= r_data[36053];
                
                r_data[36055] <= r_data[36054];
                
                r_data[36056] <= r_data[36055];
                
                r_data[36057] <= r_data[36056];
                
                r_data[36058] <= r_data[36057];
                
                r_data[36059] <= r_data[36058];
                
                r_data[36060] <= r_data[36059];
                
                r_data[36061] <= r_data[36060];
                
                r_data[36062] <= r_data[36061];
                
                r_data[36063] <= r_data[36062];
                
                r_data[36064] <= r_data[36063];
                
                r_data[36065] <= r_data[36064];
                
                r_data[36066] <= r_data[36065];
                
                r_data[36067] <= r_data[36066];
                
                r_data[36068] <= r_data[36067];
                
                r_data[36069] <= r_data[36068];
                
                r_data[36070] <= r_data[36069];
                
                r_data[36071] <= r_data[36070];
                
                r_data[36072] <= r_data[36071];
                
                r_data[36073] <= r_data[36072];
                
                r_data[36074] <= r_data[36073];
                
                r_data[36075] <= r_data[36074];
                
                r_data[36076] <= r_data[36075];
                
                r_data[36077] <= r_data[36076];
                
                r_data[36078] <= r_data[36077];
                
                r_data[36079] <= r_data[36078];
                
                r_data[36080] <= r_data[36079];
                
                r_data[36081] <= r_data[36080];
                
                r_data[36082] <= r_data[36081];
                
                r_data[36083] <= r_data[36082];
                
                r_data[36084] <= r_data[36083];
                
                r_data[36085] <= r_data[36084];
                
                r_data[36086] <= r_data[36085];
                
                r_data[36087] <= r_data[36086];
                
                r_data[36088] <= r_data[36087];
                
                r_data[36089] <= r_data[36088];
                
                r_data[36090] <= r_data[36089];
                
                r_data[36091] <= r_data[36090];
                
                r_data[36092] <= r_data[36091];
                
                r_data[36093] <= r_data[36092];
                
                r_data[36094] <= r_data[36093];
                
                r_data[36095] <= r_data[36094];
                
                r_data[36096] <= r_data[36095];
                
                r_data[36097] <= r_data[36096];
                
                r_data[36098] <= r_data[36097];
                
                r_data[36099] <= r_data[36098];
                
                r_data[36100] <= r_data[36099];
                
                r_data[36101] <= r_data[36100];
                
                r_data[36102] <= r_data[36101];
                
                r_data[36103] <= r_data[36102];
                
                r_data[36104] <= r_data[36103];
                
                r_data[36105] <= r_data[36104];
                
                r_data[36106] <= r_data[36105];
                
                r_data[36107] <= r_data[36106];
                
                r_data[36108] <= r_data[36107];
                
                r_data[36109] <= r_data[36108];
                
                r_data[36110] <= r_data[36109];
                
                r_data[36111] <= r_data[36110];
                
                r_data[36112] <= r_data[36111];
                
                r_data[36113] <= r_data[36112];
                
                r_data[36114] <= r_data[36113];
                
                r_data[36115] <= r_data[36114];
                
                r_data[36116] <= r_data[36115];
                
                r_data[36117] <= r_data[36116];
                
                r_data[36118] <= r_data[36117];
                
                r_data[36119] <= r_data[36118];
                
                r_data[36120] <= r_data[36119];
                
                r_data[36121] <= r_data[36120];
                
                r_data[36122] <= r_data[36121];
                
                r_data[36123] <= r_data[36122];
                
                r_data[36124] <= r_data[36123];
                
                r_data[36125] <= r_data[36124];
                
                r_data[36126] <= r_data[36125];
                
                r_data[36127] <= r_data[36126];
                
                r_data[36128] <= r_data[36127];
                
                r_data[36129] <= r_data[36128];
                
                r_data[36130] <= r_data[36129];
                
                r_data[36131] <= r_data[36130];
                
                r_data[36132] <= r_data[36131];
                
                r_data[36133] <= r_data[36132];
                
                r_data[36134] <= r_data[36133];
                
                r_data[36135] <= r_data[36134];
                
                r_data[36136] <= r_data[36135];
                
                r_data[36137] <= r_data[36136];
                
                r_data[36138] <= r_data[36137];
                
                r_data[36139] <= r_data[36138];
                
                r_data[36140] <= r_data[36139];
                
                r_data[36141] <= r_data[36140];
                
                r_data[36142] <= r_data[36141];
                
                r_data[36143] <= r_data[36142];
                
                r_data[36144] <= r_data[36143];
                
                r_data[36145] <= r_data[36144];
                
                r_data[36146] <= r_data[36145];
                
                r_data[36147] <= r_data[36146];
                
                r_data[36148] <= r_data[36147];
                
                r_data[36149] <= r_data[36148];
                
                r_data[36150] <= r_data[36149];
                
                r_data[36151] <= r_data[36150];
                
                r_data[36152] <= r_data[36151];
                
                r_data[36153] <= r_data[36152];
                
                r_data[36154] <= r_data[36153];
                
                r_data[36155] <= r_data[36154];
                
                r_data[36156] <= r_data[36155];
                
                r_data[36157] <= r_data[36156];
                
                r_data[36158] <= r_data[36157];
                
                r_data[36159] <= r_data[36158];
                
                r_data[36160] <= r_data[36159];
                
                r_data[36161] <= r_data[36160];
                
                r_data[36162] <= r_data[36161];
                
                r_data[36163] <= r_data[36162];
                
                r_data[36164] <= r_data[36163];
                
                r_data[36165] <= r_data[36164];
                
                r_data[36166] <= r_data[36165];
                
                r_data[36167] <= r_data[36166];
                
                r_data[36168] <= r_data[36167];
                
                r_data[36169] <= r_data[36168];
                
                r_data[36170] <= r_data[36169];
                
                r_data[36171] <= r_data[36170];
                
                r_data[36172] <= r_data[36171];
                
                r_data[36173] <= r_data[36172];
                
                r_data[36174] <= r_data[36173];
                
                r_data[36175] <= r_data[36174];
                
                r_data[36176] <= r_data[36175];
                
                r_data[36177] <= r_data[36176];
                
                r_data[36178] <= r_data[36177];
                
                r_data[36179] <= r_data[36178];
                
                r_data[36180] <= r_data[36179];
                
                r_data[36181] <= r_data[36180];
                
                r_data[36182] <= r_data[36181];
                
                r_data[36183] <= r_data[36182];
                
                r_data[36184] <= r_data[36183];
                
                r_data[36185] <= r_data[36184];
                
                r_data[36186] <= r_data[36185];
                
                r_data[36187] <= r_data[36186];
                
                r_data[36188] <= r_data[36187];
                
                r_data[36189] <= r_data[36188];
                
                r_data[36190] <= r_data[36189];
                
                r_data[36191] <= r_data[36190];
                
                r_data[36192] <= r_data[36191];
                
                r_data[36193] <= r_data[36192];
                
                r_data[36194] <= r_data[36193];
                
                r_data[36195] <= r_data[36194];
                
                r_data[36196] <= r_data[36195];
                
                r_data[36197] <= r_data[36196];
                
                r_data[36198] <= r_data[36197];
                
                r_data[36199] <= r_data[36198];
                
                r_data[36200] <= r_data[36199];
                
                r_data[36201] <= r_data[36200];
                
                r_data[36202] <= r_data[36201];
                
                r_data[36203] <= r_data[36202];
                
                r_data[36204] <= r_data[36203];
                
                r_data[36205] <= r_data[36204];
                
                r_data[36206] <= r_data[36205];
                
                r_data[36207] <= r_data[36206];
                
                r_data[36208] <= r_data[36207];
                
                r_data[36209] <= r_data[36208];
                
                r_data[36210] <= r_data[36209];
                
                r_data[36211] <= r_data[36210];
                
                r_data[36212] <= r_data[36211];
                
                r_data[36213] <= r_data[36212];
                
                r_data[36214] <= r_data[36213];
                
                r_data[36215] <= r_data[36214];
                
                r_data[36216] <= r_data[36215];
                
                r_data[36217] <= r_data[36216];
                
                r_data[36218] <= r_data[36217];
                
                r_data[36219] <= r_data[36218];
                
                r_data[36220] <= r_data[36219];
                
                r_data[36221] <= r_data[36220];
                
                r_data[36222] <= r_data[36221];
                
                r_data[36223] <= r_data[36222];
                
                r_data[36224] <= r_data[36223];
                
                r_data[36225] <= r_data[36224];
                
                r_data[36226] <= r_data[36225];
                
                r_data[36227] <= r_data[36226];
                
                r_data[36228] <= r_data[36227];
                
                r_data[36229] <= r_data[36228];
                
                r_data[36230] <= r_data[36229];
                
                r_data[36231] <= r_data[36230];
                
                r_data[36232] <= r_data[36231];
                
                r_data[36233] <= r_data[36232];
                
                r_data[36234] <= r_data[36233];
                
                r_data[36235] <= r_data[36234];
                
                r_data[36236] <= r_data[36235];
                
                r_data[36237] <= r_data[36236];
                
                r_data[36238] <= r_data[36237];
                
                r_data[36239] <= r_data[36238];
                
                r_data[36240] <= r_data[36239];
                
                r_data[36241] <= r_data[36240];
                
                r_data[36242] <= r_data[36241];
                
                r_data[36243] <= r_data[36242];
                
                r_data[36244] <= r_data[36243];
                
                r_data[36245] <= r_data[36244];
                
                r_data[36246] <= r_data[36245];
                
                r_data[36247] <= r_data[36246];
                
                r_data[36248] <= r_data[36247];
                
                r_data[36249] <= r_data[36248];
                
                r_data[36250] <= r_data[36249];
                
                r_data[36251] <= r_data[36250];
                
                r_data[36252] <= r_data[36251];
                
                r_data[36253] <= r_data[36252];
                
                r_data[36254] <= r_data[36253];
                
                r_data[36255] <= r_data[36254];
                
                r_data[36256] <= r_data[36255];
                
                r_data[36257] <= r_data[36256];
                
                r_data[36258] <= r_data[36257];
                
                r_data[36259] <= r_data[36258];
                
                r_data[36260] <= r_data[36259];
                
                r_data[36261] <= r_data[36260];
                
                r_data[36262] <= r_data[36261];
                
                r_data[36263] <= r_data[36262];
                
                r_data[36264] <= r_data[36263];
                
                r_data[36265] <= r_data[36264];
                
                r_data[36266] <= r_data[36265];
                
                r_data[36267] <= r_data[36266];
                
                r_data[36268] <= r_data[36267];
                
                r_data[36269] <= r_data[36268];
                
                r_data[36270] <= r_data[36269];
                
                r_data[36271] <= r_data[36270];
                
                r_data[36272] <= r_data[36271];
                
                r_data[36273] <= r_data[36272];
                
                r_data[36274] <= r_data[36273];
                
                r_data[36275] <= r_data[36274];
                
                r_data[36276] <= r_data[36275];
                
                r_data[36277] <= r_data[36276];
                
                r_data[36278] <= r_data[36277];
                
                r_data[36279] <= r_data[36278];
                
                r_data[36280] <= r_data[36279];
                
                r_data[36281] <= r_data[36280];
                
                r_data[36282] <= r_data[36281];
                
                r_data[36283] <= r_data[36282];
                
                r_data[36284] <= r_data[36283];
                
                r_data[36285] <= r_data[36284];
                
                r_data[36286] <= r_data[36285];
                
                r_data[36287] <= r_data[36286];
                
                r_data[36288] <= r_data[36287];
                
                r_data[36289] <= r_data[36288];
                
                r_data[36290] <= r_data[36289];
                
                r_data[36291] <= r_data[36290];
                
                r_data[36292] <= r_data[36291];
                
                r_data[36293] <= r_data[36292];
                
                r_data[36294] <= r_data[36293];
                
                r_data[36295] <= r_data[36294];
                
                r_data[36296] <= r_data[36295];
                
                r_data[36297] <= r_data[36296];
                
                r_data[36298] <= r_data[36297];
                
                r_data[36299] <= r_data[36298];
                
                r_data[36300] <= r_data[36299];
                
                r_data[36301] <= r_data[36300];
                
                r_data[36302] <= r_data[36301];
                
                r_data[36303] <= r_data[36302];
                
                r_data[36304] <= r_data[36303];
                
                r_data[36305] <= r_data[36304];
                
                r_data[36306] <= r_data[36305];
                
                r_data[36307] <= r_data[36306];
                
                r_data[36308] <= r_data[36307];
                
                r_data[36309] <= r_data[36308];
                
                r_data[36310] <= r_data[36309];
                
                r_data[36311] <= r_data[36310];
                
                r_data[36312] <= r_data[36311];
                
                r_data[36313] <= r_data[36312];
                
                r_data[36314] <= r_data[36313];
                
                r_data[36315] <= r_data[36314];
                
                r_data[36316] <= r_data[36315];
                
                r_data[36317] <= r_data[36316];
                
                r_data[36318] <= r_data[36317];
                
                r_data[36319] <= r_data[36318];
                
                r_data[36320] <= r_data[36319];
                
                r_data[36321] <= r_data[36320];
                
                r_data[36322] <= r_data[36321];
                
                r_data[36323] <= r_data[36322];
                
                r_data[36324] <= r_data[36323];
                
                r_data[36325] <= r_data[36324];
                
                r_data[36326] <= r_data[36325];
                
                r_data[36327] <= r_data[36326];
                
                r_data[36328] <= r_data[36327];
                
                r_data[36329] <= r_data[36328];
                
                r_data[36330] <= r_data[36329];
                
                r_data[36331] <= r_data[36330];
                
                r_data[36332] <= r_data[36331];
                
                r_data[36333] <= r_data[36332];
                
                r_data[36334] <= r_data[36333];
                
                r_data[36335] <= r_data[36334];
                
                r_data[36336] <= r_data[36335];
                
                r_data[36337] <= r_data[36336];
                
                r_data[36338] <= r_data[36337];
                
                r_data[36339] <= r_data[36338];
                
                r_data[36340] <= r_data[36339];
                
                r_data[36341] <= r_data[36340];
                
                r_data[36342] <= r_data[36341];
                
                r_data[36343] <= r_data[36342];
                
                r_data[36344] <= r_data[36343];
                
                r_data[36345] <= r_data[36344];
                
                r_data[36346] <= r_data[36345];
                
                r_data[36347] <= r_data[36346];
                
                r_data[36348] <= r_data[36347];
                
                r_data[36349] <= r_data[36348];
                
                r_data[36350] <= r_data[36349];
                
                r_data[36351] <= r_data[36350];
                
                r_data[36352] <= r_data[36351];
                
                r_data[36353] <= r_data[36352];
                
                r_data[36354] <= r_data[36353];
                
                r_data[36355] <= r_data[36354];
                
                r_data[36356] <= r_data[36355];
                
                r_data[36357] <= r_data[36356];
                
                r_data[36358] <= r_data[36357];
                
                r_data[36359] <= r_data[36358];
                
                r_data[36360] <= r_data[36359];
                
                r_data[36361] <= r_data[36360];
                
                r_data[36362] <= r_data[36361];
                
                r_data[36363] <= r_data[36362];
                
                r_data[36364] <= r_data[36363];
                
                r_data[36365] <= r_data[36364];
                
                r_data[36366] <= r_data[36365];
                
                r_data[36367] <= r_data[36366];
                
                r_data[36368] <= r_data[36367];
                
                r_data[36369] <= r_data[36368];
                
                r_data[36370] <= r_data[36369];
                
                r_data[36371] <= r_data[36370];
                
                r_data[36372] <= r_data[36371];
                
                r_data[36373] <= r_data[36372];
                
                r_data[36374] <= r_data[36373];
                
                r_data[36375] <= r_data[36374];
                
                r_data[36376] <= r_data[36375];
                
                r_data[36377] <= r_data[36376];
                
                r_data[36378] <= r_data[36377];
                
                r_data[36379] <= r_data[36378];
                
                r_data[36380] <= r_data[36379];
                
                r_data[36381] <= r_data[36380];
                
                r_data[36382] <= r_data[36381];
                
                r_data[36383] <= r_data[36382];
                
                r_data[36384] <= r_data[36383];
                
                r_data[36385] <= r_data[36384];
                
                r_data[36386] <= r_data[36385];
                
                r_data[36387] <= r_data[36386];
                
                r_data[36388] <= r_data[36387];
                
                r_data[36389] <= r_data[36388];
                
                r_data[36390] <= r_data[36389];
                
                r_data[36391] <= r_data[36390];
                
                r_data[36392] <= r_data[36391];
                
                r_data[36393] <= r_data[36392];
                
                r_data[36394] <= r_data[36393];
                
                r_data[36395] <= r_data[36394];
                
                r_data[36396] <= r_data[36395];
                
                r_data[36397] <= r_data[36396];
                
                r_data[36398] <= r_data[36397];
                
                r_data[36399] <= r_data[36398];
                
                r_data[36400] <= r_data[36399];
                
                r_data[36401] <= r_data[36400];
                
                r_data[36402] <= r_data[36401];
                
                r_data[36403] <= r_data[36402];
                
                r_data[36404] <= r_data[36403];
                
                r_data[36405] <= r_data[36404];
                
                r_data[36406] <= r_data[36405];
                
                r_data[36407] <= r_data[36406];
                
                r_data[36408] <= r_data[36407];
                
                r_data[36409] <= r_data[36408];
                
                r_data[36410] <= r_data[36409];
                
                r_data[36411] <= r_data[36410];
                
                r_data[36412] <= r_data[36411];
                
                r_data[36413] <= r_data[36412];
                
                r_data[36414] <= r_data[36413];
                
                r_data[36415] <= r_data[36414];
                
                r_data[36416] <= r_data[36415];
                
                r_data[36417] <= r_data[36416];
                
                r_data[36418] <= r_data[36417];
                
                r_data[36419] <= r_data[36418];
                
                r_data[36420] <= r_data[36419];
                
                r_data[36421] <= r_data[36420];
                
                r_data[36422] <= r_data[36421];
                
                r_data[36423] <= r_data[36422];
                
                r_data[36424] <= r_data[36423];
                
                r_data[36425] <= r_data[36424];
                
                r_data[36426] <= r_data[36425];
                
                r_data[36427] <= r_data[36426];
                
                r_data[36428] <= r_data[36427];
                
                r_data[36429] <= r_data[36428];
                
                r_data[36430] <= r_data[36429];
                
                r_data[36431] <= r_data[36430];
                
                r_data[36432] <= r_data[36431];
                
                r_data[36433] <= r_data[36432];
                
                r_data[36434] <= r_data[36433];
                
                r_data[36435] <= r_data[36434];
                
                r_data[36436] <= r_data[36435];
                
                r_data[36437] <= r_data[36436];
                
                r_data[36438] <= r_data[36437];
                
                r_data[36439] <= r_data[36438];
                
                r_data[36440] <= r_data[36439];
                
                r_data[36441] <= r_data[36440];
                
                r_data[36442] <= r_data[36441];
                
                r_data[36443] <= r_data[36442];
                
                r_data[36444] <= r_data[36443];
                
                r_data[36445] <= r_data[36444];
                
                r_data[36446] <= r_data[36445];
                
                r_data[36447] <= r_data[36446];
                
                r_data[36448] <= r_data[36447];
                
                r_data[36449] <= r_data[36448];
                
                r_data[36450] <= r_data[36449];
                
                r_data[36451] <= r_data[36450];
                
                r_data[36452] <= r_data[36451];
                
                r_data[36453] <= r_data[36452];
                
                r_data[36454] <= r_data[36453];
                
                r_data[36455] <= r_data[36454];
                
                r_data[36456] <= r_data[36455];
                
                r_data[36457] <= r_data[36456];
                
                r_data[36458] <= r_data[36457];
                
                r_data[36459] <= r_data[36458];
                
                r_data[36460] <= r_data[36459];
                
                r_data[36461] <= r_data[36460];
                
                r_data[36462] <= r_data[36461];
                
                r_data[36463] <= r_data[36462];
                
                r_data[36464] <= r_data[36463];
                
                r_data[36465] <= r_data[36464];
                
                r_data[36466] <= r_data[36465];
                
                r_data[36467] <= r_data[36466];
                
                r_data[36468] <= r_data[36467];
                
                r_data[36469] <= r_data[36468];
                
                r_data[36470] <= r_data[36469];
                
                r_data[36471] <= r_data[36470];
                
                r_data[36472] <= r_data[36471];
                
                r_data[36473] <= r_data[36472];
                
                r_data[36474] <= r_data[36473];
                
                r_data[36475] <= r_data[36474];
                
                r_data[36476] <= r_data[36475];
                
                r_data[36477] <= r_data[36476];
                
                r_data[36478] <= r_data[36477];
                
                r_data[36479] <= r_data[36478];
                
                r_data[36480] <= r_data[36479];
                
                r_data[36481] <= r_data[36480];
                
                r_data[36482] <= r_data[36481];
                
                r_data[36483] <= r_data[36482];
                
                r_data[36484] <= r_data[36483];
                
                r_data[36485] <= r_data[36484];
                
                r_data[36486] <= r_data[36485];
                
                r_data[36487] <= r_data[36486];
                
                r_data[36488] <= r_data[36487];
                
                r_data[36489] <= r_data[36488];
                
                r_data[36490] <= r_data[36489];
                
                r_data[36491] <= r_data[36490];
                
                r_data[36492] <= r_data[36491];
                
                r_data[36493] <= r_data[36492];
                
                r_data[36494] <= r_data[36493];
                
                r_data[36495] <= r_data[36494];
                
                r_data[36496] <= r_data[36495];
                
                r_data[36497] <= r_data[36496];
                
                r_data[36498] <= r_data[36497];
                
                r_data[36499] <= r_data[36498];
                
                r_data[36500] <= r_data[36499];
                
                r_data[36501] <= r_data[36500];
                
                r_data[36502] <= r_data[36501];
                
                r_data[36503] <= r_data[36502];
                
                r_data[36504] <= r_data[36503];
                
                r_data[36505] <= r_data[36504];
                
                r_data[36506] <= r_data[36505];
                
                r_data[36507] <= r_data[36506];
                
                r_data[36508] <= r_data[36507];
                
                r_data[36509] <= r_data[36508];
                
                r_data[36510] <= r_data[36509];
                
                r_data[36511] <= r_data[36510];
                
                r_data[36512] <= r_data[36511];
                
                r_data[36513] <= r_data[36512];
                
                r_data[36514] <= r_data[36513];
                
                r_data[36515] <= r_data[36514];
                
                r_data[36516] <= r_data[36515];
                
                r_data[36517] <= r_data[36516];
                
                r_data[36518] <= r_data[36517];
                
                r_data[36519] <= r_data[36518];
                
                r_data[36520] <= r_data[36519];
                
                r_data[36521] <= r_data[36520];
                
                r_data[36522] <= r_data[36521];
                
                r_data[36523] <= r_data[36522];
                
                r_data[36524] <= r_data[36523];
                
                r_data[36525] <= r_data[36524];
                
                r_data[36526] <= r_data[36525];
                
                r_data[36527] <= r_data[36526];
                
                r_data[36528] <= r_data[36527];
                
                r_data[36529] <= r_data[36528];
                
                r_data[36530] <= r_data[36529];
                
                r_data[36531] <= r_data[36530];
                
                r_data[36532] <= r_data[36531];
                
                r_data[36533] <= r_data[36532];
                
                r_data[36534] <= r_data[36533];
                
                r_data[36535] <= r_data[36534];
                
                r_data[36536] <= r_data[36535];
                
                r_data[36537] <= r_data[36536];
                
                r_data[36538] <= r_data[36537];
                
                r_data[36539] <= r_data[36538];
                
                r_data[36540] <= r_data[36539];
                
                r_data[36541] <= r_data[36540];
                
                r_data[36542] <= r_data[36541];
                
                r_data[36543] <= r_data[36542];
                
                r_data[36544] <= r_data[36543];
                
                r_data[36545] <= r_data[36544];
                
                r_data[36546] <= r_data[36545];
                
                r_data[36547] <= r_data[36546];
                
                r_data[36548] <= r_data[36547];
                
                r_data[36549] <= r_data[36548];
                
                r_data[36550] <= r_data[36549];
                
                r_data[36551] <= r_data[36550];
                
                r_data[36552] <= r_data[36551];
                
                r_data[36553] <= r_data[36552];
                
                r_data[36554] <= r_data[36553];
                
                r_data[36555] <= r_data[36554];
                
                r_data[36556] <= r_data[36555];
                
                r_data[36557] <= r_data[36556];
                
                r_data[36558] <= r_data[36557];
                
                r_data[36559] <= r_data[36558];
                
                r_data[36560] <= r_data[36559];
                
                r_data[36561] <= r_data[36560];
                
                r_data[36562] <= r_data[36561];
                
                r_data[36563] <= r_data[36562];
                
                r_data[36564] <= r_data[36563];
                
                r_data[36565] <= r_data[36564];
                
                r_data[36566] <= r_data[36565];
                
                r_data[36567] <= r_data[36566];
                
                r_data[36568] <= r_data[36567];
                
                r_data[36569] <= r_data[36568];
                
                r_data[36570] <= r_data[36569];
                
                r_data[36571] <= r_data[36570];
                
                r_data[36572] <= r_data[36571];
                
                r_data[36573] <= r_data[36572];
                
                r_data[36574] <= r_data[36573];
                
                r_data[36575] <= r_data[36574];
                
                r_data[36576] <= r_data[36575];
                
                r_data[36577] <= r_data[36576];
                
                r_data[36578] <= r_data[36577];
                
                r_data[36579] <= r_data[36578];
                
                r_data[36580] <= r_data[36579];
                
                r_data[36581] <= r_data[36580];
                
                r_data[36582] <= r_data[36581];
                
                r_data[36583] <= r_data[36582];
                
                r_data[36584] <= r_data[36583];
                
                r_data[36585] <= r_data[36584];
                
                r_data[36586] <= r_data[36585];
                
                r_data[36587] <= r_data[36586];
                
                r_data[36588] <= r_data[36587];
                
                r_data[36589] <= r_data[36588];
                
                r_data[36590] <= r_data[36589];
                
                r_data[36591] <= r_data[36590];
                
                r_data[36592] <= r_data[36591];
                
                r_data[36593] <= r_data[36592];
                
                r_data[36594] <= r_data[36593];
                
                r_data[36595] <= r_data[36594];
                
                r_data[36596] <= r_data[36595];
                
                r_data[36597] <= r_data[36596];
                
                r_data[36598] <= r_data[36597];
                
                r_data[36599] <= r_data[36598];
                
                r_data[36600] <= r_data[36599];
                
                r_data[36601] <= r_data[36600];
                
                r_data[36602] <= r_data[36601];
                
                r_data[36603] <= r_data[36602];
                
                r_data[36604] <= r_data[36603];
                
                r_data[36605] <= r_data[36604];
                
                r_data[36606] <= r_data[36605];
                
                r_data[36607] <= r_data[36606];
                
                r_data[36608] <= r_data[36607];
                
                r_data[36609] <= r_data[36608];
                
                r_data[36610] <= r_data[36609];
                
                r_data[36611] <= r_data[36610];
                
                r_data[36612] <= r_data[36611];
                
                r_data[36613] <= r_data[36612];
                
                r_data[36614] <= r_data[36613];
                
                r_data[36615] <= r_data[36614];
                
                r_data[36616] <= r_data[36615];
                
                r_data[36617] <= r_data[36616];
                
                r_data[36618] <= r_data[36617];
                
                r_data[36619] <= r_data[36618];
                
                r_data[36620] <= r_data[36619];
                
                r_data[36621] <= r_data[36620];
                
                r_data[36622] <= r_data[36621];
                
                r_data[36623] <= r_data[36622];
                
                r_data[36624] <= r_data[36623];
                
                r_data[36625] <= r_data[36624];
                
                r_data[36626] <= r_data[36625];
                
                r_data[36627] <= r_data[36626];
                
                r_data[36628] <= r_data[36627];
                
                r_data[36629] <= r_data[36628];
                
                r_data[36630] <= r_data[36629];
                
                r_data[36631] <= r_data[36630];
                
                r_data[36632] <= r_data[36631];
                
                r_data[36633] <= r_data[36632];
                
                r_data[36634] <= r_data[36633];
                
                r_data[36635] <= r_data[36634];
                
                r_data[36636] <= r_data[36635];
                
                r_data[36637] <= r_data[36636];
                
                r_data[36638] <= r_data[36637];
                
                r_data[36639] <= r_data[36638];
                
                r_data[36640] <= r_data[36639];
                
                r_data[36641] <= r_data[36640];
                
                r_data[36642] <= r_data[36641];
                
                r_data[36643] <= r_data[36642];
                
                r_data[36644] <= r_data[36643];
                
                r_data[36645] <= r_data[36644];
                
                r_data[36646] <= r_data[36645];
                
                r_data[36647] <= r_data[36646];
                
                r_data[36648] <= r_data[36647];
                
                r_data[36649] <= r_data[36648];
                
                r_data[36650] <= r_data[36649];
                
                r_data[36651] <= r_data[36650];
                
                r_data[36652] <= r_data[36651];
                
                r_data[36653] <= r_data[36652];
                
                r_data[36654] <= r_data[36653];
                
                r_data[36655] <= r_data[36654];
                
                r_data[36656] <= r_data[36655];
                
                r_data[36657] <= r_data[36656];
                
                r_data[36658] <= r_data[36657];
                
                r_data[36659] <= r_data[36658];
                
                r_data[36660] <= r_data[36659];
                
                r_data[36661] <= r_data[36660];
                
                r_data[36662] <= r_data[36661];
                
                r_data[36663] <= r_data[36662];
                
                r_data[36664] <= r_data[36663];
                
                r_data[36665] <= r_data[36664];
                
                r_data[36666] <= r_data[36665];
                
                r_data[36667] <= r_data[36666];
                
                r_data[36668] <= r_data[36667];
                
                r_data[36669] <= r_data[36668];
                
                r_data[36670] <= r_data[36669];
                
                r_data[36671] <= r_data[36670];
                
                r_data[36672] <= r_data[36671];
                
                r_data[36673] <= r_data[36672];
                
                r_data[36674] <= r_data[36673];
                
                r_data[36675] <= r_data[36674];
                
                r_data[36676] <= r_data[36675];
                
                r_data[36677] <= r_data[36676];
                
                r_data[36678] <= r_data[36677];
                
                r_data[36679] <= r_data[36678];
                
                r_data[36680] <= r_data[36679];
                
                r_data[36681] <= r_data[36680];
                
                r_data[36682] <= r_data[36681];
                
                r_data[36683] <= r_data[36682];
                
                r_data[36684] <= r_data[36683];
                
                r_data[36685] <= r_data[36684];
                
                r_data[36686] <= r_data[36685];
                
                r_data[36687] <= r_data[36686];
                
                r_data[36688] <= r_data[36687];
                
                r_data[36689] <= r_data[36688];
                
                r_data[36690] <= r_data[36689];
                
                r_data[36691] <= r_data[36690];
                
                r_data[36692] <= r_data[36691];
                
                r_data[36693] <= r_data[36692];
                
                r_data[36694] <= r_data[36693];
                
                r_data[36695] <= r_data[36694];
                
                r_data[36696] <= r_data[36695];
                
                r_data[36697] <= r_data[36696];
                
                r_data[36698] <= r_data[36697];
                
                r_data[36699] <= r_data[36698];
                
                r_data[36700] <= r_data[36699];
                
                r_data[36701] <= r_data[36700];
                
                r_data[36702] <= r_data[36701];
                
                r_data[36703] <= r_data[36702];
                
                r_data[36704] <= r_data[36703];
                
                r_data[36705] <= r_data[36704];
                
                r_data[36706] <= r_data[36705];
                
                r_data[36707] <= r_data[36706];
                
                r_data[36708] <= r_data[36707];
                
                r_data[36709] <= r_data[36708];
                
                r_data[36710] <= r_data[36709];
                
                r_data[36711] <= r_data[36710];
                
                r_data[36712] <= r_data[36711];
                
                r_data[36713] <= r_data[36712];
                
                r_data[36714] <= r_data[36713];
                
                r_data[36715] <= r_data[36714];
                
                r_data[36716] <= r_data[36715];
                
                r_data[36717] <= r_data[36716];
                
                r_data[36718] <= r_data[36717];
                
                r_data[36719] <= r_data[36718];
                
                r_data[36720] <= r_data[36719];
                
                r_data[36721] <= r_data[36720];
                
                r_data[36722] <= r_data[36721];
                
                r_data[36723] <= r_data[36722];
                
                r_data[36724] <= r_data[36723];
                
                r_data[36725] <= r_data[36724];
                
                r_data[36726] <= r_data[36725];
                
                r_data[36727] <= r_data[36726];
                
                r_data[36728] <= r_data[36727];
                
                r_data[36729] <= r_data[36728];
                
                r_data[36730] <= r_data[36729];
                
                r_data[36731] <= r_data[36730];
                
                r_data[36732] <= r_data[36731];
                
                r_data[36733] <= r_data[36732];
                
                r_data[36734] <= r_data[36733];
                
                r_data[36735] <= r_data[36734];
                
                r_data[36736] <= r_data[36735];
                
                r_data[36737] <= r_data[36736];
                
                r_data[36738] <= r_data[36737];
                
                r_data[36739] <= r_data[36738];
                
                r_data[36740] <= r_data[36739];
                
                r_data[36741] <= r_data[36740];
                
                r_data[36742] <= r_data[36741];
                
                r_data[36743] <= r_data[36742];
                
                r_data[36744] <= r_data[36743];
                
                r_data[36745] <= r_data[36744];
                
                r_data[36746] <= r_data[36745];
                
                r_data[36747] <= r_data[36746];
                
                r_data[36748] <= r_data[36747];
                
                r_data[36749] <= r_data[36748];
                
                r_data[36750] <= r_data[36749];
                
                r_data[36751] <= r_data[36750];
                
                r_data[36752] <= r_data[36751];
                
                r_data[36753] <= r_data[36752];
                
                r_data[36754] <= r_data[36753];
                
                r_data[36755] <= r_data[36754];
                
                r_data[36756] <= r_data[36755];
                
                r_data[36757] <= r_data[36756];
                
                r_data[36758] <= r_data[36757];
                
                r_data[36759] <= r_data[36758];
                
                r_data[36760] <= r_data[36759];
                
                r_data[36761] <= r_data[36760];
                
                r_data[36762] <= r_data[36761];
                
                r_data[36763] <= r_data[36762];
                
                r_data[36764] <= r_data[36763];
                
                r_data[36765] <= r_data[36764];
                
                r_data[36766] <= r_data[36765];
                
                r_data[36767] <= r_data[36766];
                
                r_data[36768] <= r_data[36767];
                
                r_data[36769] <= r_data[36768];
                
                r_data[36770] <= r_data[36769];
                
                r_data[36771] <= r_data[36770];
                
                r_data[36772] <= r_data[36771];
                
                r_data[36773] <= r_data[36772];
                
                r_data[36774] <= r_data[36773];
                
                r_data[36775] <= r_data[36774];
                
                r_data[36776] <= r_data[36775];
                
                r_data[36777] <= r_data[36776];
                
                r_data[36778] <= r_data[36777];
                
                r_data[36779] <= r_data[36778];
                
                r_data[36780] <= r_data[36779];
                
                r_data[36781] <= r_data[36780];
                
                r_data[36782] <= r_data[36781];
                
                r_data[36783] <= r_data[36782];
                
                r_data[36784] <= r_data[36783];
                
                r_data[36785] <= r_data[36784];
                
                r_data[36786] <= r_data[36785];
                
                r_data[36787] <= r_data[36786];
                
                r_data[36788] <= r_data[36787];
                
                r_data[36789] <= r_data[36788];
                
                r_data[36790] <= r_data[36789];
                
                r_data[36791] <= r_data[36790];
                
                r_data[36792] <= r_data[36791];
                
                r_data[36793] <= r_data[36792];
                
                r_data[36794] <= r_data[36793];
                
                r_data[36795] <= r_data[36794];
                
                r_data[36796] <= r_data[36795];
                
                r_data[36797] <= r_data[36796];
                
                r_data[36798] <= r_data[36797];
                
                r_data[36799] <= r_data[36798];
                
                r_data[36800] <= r_data[36799];
                
                r_data[36801] <= r_data[36800];
                
                r_data[36802] <= r_data[36801];
                
                r_data[36803] <= r_data[36802];
                
                r_data[36804] <= r_data[36803];
                
                r_data[36805] <= r_data[36804];
                
                r_data[36806] <= r_data[36805];
                
                r_data[36807] <= r_data[36806];
                
                r_data[36808] <= r_data[36807];
                
                r_data[36809] <= r_data[36808];
                
                r_data[36810] <= r_data[36809];
                
                r_data[36811] <= r_data[36810];
                
                r_data[36812] <= r_data[36811];
                
                r_data[36813] <= r_data[36812];
                
                r_data[36814] <= r_data[36813];
                
                r_data[36815] <= r_data[36814];
                
                r_data[36816] <= r_data[36815];
                
                r_data[36817] <= r_data[36816];
                
                r_data[36818] <= r_data[36817];
                
                r_data[36819] <= r_data[36818];
                
                r_data[36820] <= r_data[36819];
                
                r_data[36821] <= r_data[36820];
                
                r_data[36822] <= r_data[36821];
                
                r_data[36823] <= r_data[36822];
                
                r_data[36824] <= r_data[36823];
                
                r_data[36825] <= r_data[36824];
                
                r_data[36826] <= r_data[36825];
                
                r_data[36827] <= r_data[36826];
                
                r_data[36828] <= r_data[36827];
                
                r_data[36829] <= r_data[36828];
                
                r_data[36830] <= r_data[36829];
                
                r_data[36831] <= r_data[36830];
                
                r_data[36832] <= r_data[36831];
                
                r_data[36833] <= r_data[36832];
                
                r_data[36834] <= r_data[36833];
                
                r_data[36835] <= r_data[36834];
                
                r_data[36836] <= r_data[36835];
                
                r_data[36837] <= r_data[36836];
                
                r_data[36838] <= r_data[36837];
                
                r_data[36839] <= r_data[36838];
                
                r_data[36840] <= r_data[36839];
                
                r_data[36841] <= r_data[36840];
                
                r_data[36842] <= r_data[36841];
                
                r_data[36843] <= r_data[36842];
                
                r_data[36844] <= r_data[36843];
                
                r_data[36845] <= r_data[36844];
                
                r_data[36846] <= r_data[36845];
                
                r_data[36847] <= r_data[36846];
                
                r_data[36848] <= r_data[36847];
                
                r_data[36849] <= r_data[36848];
                
                r_data[36850] <= r_data[36849];
                
                r_data[36851] <= r_data[36850];
                
                r_data[36852] <= r_data[36851];
                
                r_data[36853] <= r_data[36852];
                
                r_data[36854] <= r_data[36853];
                
                r_data[36855] <= r_data[36854];
                
                r_data[36856] <= r_data[36855];
                
                r_data[36857] <= r_data[36856];
                
                r_data[36858] <= r_data[36857];
                
                r_data[36859] <= r_data[36858];
                
                r_data[36860] <= r_data[36859];
                
                r_data[36861] <= r_data[36860];
                
                r_data[36862] <= r_data[36861];
                
                r_data[36863] <= r_data[36862];
                
                r_data[36864] <= r_data[36863];
                
                r_data[36865] <= r_data[36864];
                
                r_data[36866] <= r_data[36865];
                
                r_data[36867] <= r_data[36866];
                
                r_data[36868] <= r_data[36867];
                
                r_data[36869] <= r_data[36868];
                
                r_data[36870] <= r_data[36869];
                
                r_data[36871] <= r_data[36870];
                
                r_data[36872] <= r_data[36871];
                
                r_data[36873] <= r_data[36872];
                
                r_data[36874] <= r_data[36873];
                
                r_data[36875] <= r_data[36874];
                
                r_data[36876] <= r_data[36875];
                
                r_data[36877] <= r_data[36876];
                
                r_data[36878] <= r_data[36877];
                
                r_data[36879] <= r_data[36878];
                
                r_data[36880] <= r_data[36879];
                
                r_data[36881] <= r_data[36880];
                
                r_data[36882] <= r_data[36881];
                
                r_data[36883] <= r_data[36882];
                
                r_data[36884] <= r_data[36883];
                
                r_data[36885] <= r_data[36884];
                
                r_data[36886] <= r_data[36885];
                
                r_data[36887] <= r_data[36886];
                
                r_data[36888] <= r_data[36887];
                
                r_data[36889] <= r_data[36888];
                
                r_data[36890] <= r_data[36889];
                
                r_data[36891] <= r_data[36890];
                
                r_data[36892] <= r_data[36891];
                
                r_data[36893] <= r_data[36892];
                
                r_data[36894] <= r_data[36893];
                
                r_data[36895] <= r_data[36894];
                
                r_data[36896] <= r_data[36895];
                
                r_data[36897] <= r_data[36896];
                
                r_data[36898] <= r_data[36897];
                
                r_data[36899] <= r_data[36898];
                
                r_data[36900] <= r_data[36899];
                
                r_data[36901] <= r_data[36900];
                
                r_data[36902] <= r_data[36901];
                
                r_data[36903] <= r_data[36902];
                
                r_data[36904] <= r_data[36903];
                
                r_data[36905] <= r_data[36904];
                
                r_data[36906] <= r_data[36905];
                
                r_data[36907] <= r_data[36906];
                
                r_data[36908] <= r_data[36907];
                
                r_data[36909] <= r_data[36908];
                
                r_data[36910] <= r_data[36909];
                
                r_data[36911] <= r_data[36910];
                
                r_data[36912] <= r_data[36911];
                
                r_data[36913] <= r_data[36912];
                
                r_data[36914] <= r_data[36913];
                
                r_data[36915] <= r_data[36914];
                
                r_data[36916] <= r_data[36915];
                
                r_data[36917] <= r_data[36916];
                
                r_data[36918] <= r_data[36917];
                
                r_data[36919] <= r_data[36918];
                
                r_data[36920] <= r_data[36919];
                
                r_data[36921] <= r_data[36920];
                
                r_data[36922] <= r_data[36921];
                
                r_data[36923] <= r_data[36922];
                
                r_data[36924] <= r_data[36923];
                
                r_data[36925] <= r_data[36924];
                
                r_data[36926] <= r_data[36925];
                
                r_data[36927] <= r_data[36926];
                
                r_data[36928] <= r_data[36927];
                
                r_data[36929] <= r_data[36928];
                
                r_data[36930] <= r_data[36929];
                
                r_data[36931] <= r_data[36930];
                
                r_data[36932] <= r_data[36931];
                
                r_data[36933] <= r_data[36932];
                
                r_data[36934] <= r_data[36933];
                
                r_data[36935] <= r_data[36934];
                
                r_data[36936] <= r_data[36935];
                
                r_data[36937] <= r_data[36936];
                
                r_data[36938] <= r_data[36937];
                
                r_data[36939] <= r_data[36938];
                
                r_data[36940] <= r_data[36939];
                
                r_data[36941] <= r_data[36940];
                
                r_data[36942] <= r_data[36941];
                
                r_data[36943] <= r_data[36942];
                
                r_data[36944] <= r_data[36943];
                
                r_data[36945] <= r_data[36944];
                
                r_data[36946] <= r_data[36945];
                
                r_data[36947] <= r_data[36946];
                
                r_data[36948] <= r_data[36947];
                
                r_data[36949] <= r_data[36948];
                
                r_data[36950] <= r_data[36949];
                
                r_data[36951] <= r_data[36950];
                
                r_data[36952] <= r_data[36951];
                
                r_data[36953] <= r_data[36952];
                
                r_data[36954] <= r_data[36953];
                
                r_data[36955] <= r_data[36954];
                
                r_data[36956] <= r_data[36955];
                
                r_data[36957] <= r_data[36956];
                
                r_data[36958] <= r_data[36957];
                
                r_data[36959] <= r_data[36958];
                
                r_data[36960] <= r_data[36959];
                
                r_data[36961] <= r_data[36960];
                
                r_data[36962] <= r_data[36961];
                
                r_data[36963] <= r_data[36962];
                
                r_data[36964] <= r_data[36963];
                
                r_data[36965] <= r_data[36964];
                
                r_data[36966] <= r_data[36965];
                
                r_data[36967] <= r_data[36966];
                
                r_data[36968] <= r_data[36967];
                
                r_data[36969] <= r_data[36968];
                
                r_data[36970] <= r_data[36969];
                
                r_data[36971] <= r_data[36970];
                
                r_data[36972] <= r_data[36971];
                
                r_data[36973] <= r_data[36972];
                
                r_data[36974] <= r_data[36973];
                
                r_data[36975] <= r_data[36974];
                
                r_data[36976] <= r_data[36975];
                
                r_data[36977] <= r_data[36976];
                
                r_data[36978] <= r_data[36977];
                
                r_data[36979] <= r_data[36978];
                
                r_data[36980] <= r_data[36979];
                
                r_data[36981] <= r_data[36980];
                
                r_data[36982] <= r_data[36981];
                
                r_data[36983] <= r_data[36982];
                
                r_data[36984] <= r_data[36983];
                
                r_data[36985] <= r_data[36984];
                
                r_data[36986] <= r_data[36985];
                
                r_data[36987] <= r_data[36986];
                
                r_data[36988] <= r_data[36987];
                
                r_data[36989] <= r_data[36988];
                
                r_data[36990] <= r_data[36989];
                
                r_data[36991] <= r_data[36990];
                
                r_data[36992] <= r_data[36991];
                
                r_data[36993] <= r_data[36992];
                
                r_data[36994] <= r_data[36993];
                
                r_data[36995] <= r_data[36994];
                
                r_data[36996] <= r_data[36995];
                
                r_data[36997] <= r_data[36996];
                
                r_data[36998] <= r_data[36997];
                
                r_data[36999] <= r_data[36998];
                
                r_data[37000] <= r_data[36999];
                
                r_data[37001] <= r_data[37000];
                
                r_data[37002] <= r_data[37001];
                
                r_data[37003] <= r_data[37002];
                
                r_data[37004] <= r_data[37003];
                
                r_data[37005] <= r_data[37004];
                
                r_data[37006] <= r_data[37005];
                
                r_data[37007] <= r_data[37006];
                
                r_data[37008] <= r_data[37007];
                
                r_data[37009] <= r_data[37008];
                
                r_data[37010] <= r_data[37009];
                
                r_data[37011] <= r_data[37010];
                
                r_data[37012] <= r_data[37011];
                
                r_data[37013] <= r_data[37012];
                
                r_data[37014] <= r_data[37013];
                
                r_data[37015] <= r_data[37014];
                
                r_data[37016] <= r_data[37015];
                
                r_data[37017] <= r_data[37016];
                
                r_data[37018] <= r_data[37017];
                
                r_data[37019] <= r_data[37018];
                
                r_data[37020] <= r_data[37019];
                
                r_data[37021] <= r_data[37020];
                
                r_data[37022] <= r_data[37021];
                
                r_data[37023] <= r_data[37022];
                
                r_data[37024] <= r_data[37023];
                
                r_data[37025] <= r_data[37024];
                
                r_data[37026] <= r_data[37025];
                
                r_data[37027] <= r_data[37026];
                
                r_data[37028] <= r_data[37027];
                
                r_data[37029] <= r_data[37028];
                
                r_data[37030] <= r_data[37029];
                
                r_data[37031] <= r_data[37030];
                
                r_data[37032] <= r_data[37031];
                
                r_data[37033] <= r_data[37032];
                
                r_data[37034] <= r_data[37033];
                
                r_data[37035] <= r_data[37034];
                
                r_data[37036] <= r_data[37035];
                
                r_data[37037] <= r_data[37036];
                
                r_data[37038] <= r_data[37037];
                
                r_data[37039] <= r_data[37038];
                
                r_data[37040] <= r_data[37039];
                
                r_data[37041] <= r_data[37040];
                
                r_data[37042] <= r_data[37041];
                
                r_data[37043] <= r_data[37042];
                
                r_data[37044] <= r_data[37043];
                
                r_data[37045] <= r_data[37044];
                
                r_data[37046] <= r_data[37045];
                
                r_data[37047] <= r_data[37046];
                
                r_data[37048] <= r_data[37047];
                
                r_data[37049] <= r_data[37048];
                
                r_data[37050] <= r_data[37049];
                
                r_data[37051] <= r_data[37050];
                
                r_data[37052] <= r_data[37051];
                
                r_data[37053] <= r_data[37052];
                
                r_data[37054] <= r_data[37053];
                
                r_data[37055] <= r_data[37054];
                
                r_data[37056] <= r_data[37055];
                
                r_data[37057] <= r_data[37056];
                
                r_data[37058] <= r_data[37057];
                
                r_data[37059] <= r_data[37058];
                
                r_data[37060] <= r_data[37059];
                
                r_data[37061] <= r_data[37060];
                
                r_data[37062] <= r_data[37061];
                
                r_data[37063] <= r_data[37062];
                
                r_data[37064] <= r_data[37063];
                
                r_data[37065] <= r_data[37064];
                
                r_data[37066] <= r_data[37065];
                
                r_data[37067] <= r_data[37066];
                
                r_data[37068] <= r_data[37067];
                
                r_data[37069] <= r_data[37068];
                
                r_data[37070] <= r_data[37069];
                
                r_data[37071] <= r_data[37070];
                
                r_data[37072] <= r_data[37071];
                
                r_data[37073] <= r_data[37072];
                
                r_data[37074] <= r_data[37073];
                
                r_data[37075] <= r_data[37074];
                
                r_data[37076] <= r_data[37075];
                
                r_data[37077] <= r_data[37076];
                
                r_data[37078] <= r_data[37077];
                
                r_data[37079] <= r_data[37078];
                
                r_data[37080] <= r_data[37079];
                
                r_data[37081] <= r_data[37080];
                
                r_data[37082] <= r_data[37081];
                
                r_data[37083] <= r_data[37082];
                
                r_data[37084] <= r_data[37083];
                
                r_data[37085] <= r_data[37084];
                
                r_data[37086] <= r_data[37085];
                
                r_data[37087] <= r_data[37086];
                
                r_data[37088] <= r_data[37087];
                
                r_data[37089] <= r_data[37088];
                
                r_data[37090] <= r_data[37089];
                
                r_data[37091] <= r_data[37090];
                
                r_data[37092] <= r_data[37091];
                
                r_data[37093] <= r_data[37092];
                
                r_data[37094] <= r_data[37093];
                
                r_data[37095] <= r_data[37094];
                
                r_data[37096] <= r_data[37095];
                
                r_data[37097] <= r_data[37096];
                
                r_data[37098] <= r_data[37097];
                
                r_data[37099] <= r_data[37098];
                
                r_data[37100] <= r_data[37099];
                
                r_data[37101] <= r_data[37100];
                
                r_data[37102] <= r_data[37101];
                
                r_data[37103] <= r_data[37102];
                
                r_data[37104] <= r_data[37103];
                
                r_data[37105] <= r_data[37104];
                
                r_data[37106] <= r_data[37105];
                
                r_data[37107] <= r_data[37106];
                
                r_data[37108] <= r_data[37107];
                
                r_data[37109] <= r_data[37108];
                
                r_data[37110] <= r_data[37109];
                
                r_data[37111] <= r_data[37110];
                
                r_data[37112] <= r_data[37111];
                
                r_data[37113] <= r_data[37112];
                
                r_data[37114] <= r_data[37113];
                
                r_data[37115] <= r_data[37114];
                
                r_data[37116] <= r_data[37115];
                
                r_data[37117] <= r_data[37116];
                
                r_data[37118] <= r_data[37117];
                
                r_data[37119] <= r_data[37118];
                
                r_data[37120] <= r_data[37119];
                
                r_data[37121] <= r_data[37120];
                
                r_data[37122] <= r_data[37121];
                
                r_data[37123] <= r_data[37122];
                
                r_data[37124] <= r_data[37123];
                
                r_data[37125] <= r_data[37124];
                
                r_data[37126] <= r_data[37125];
                
                r_data[37127] <= r_data[37126];
                
                r_data[37128] <= r_data[37127];
                
                r_data[37129] <= r_data[37128];
                
                r_data[37130] <= r_data[37129];
                
                r_data[37131] <= r_data[37130];
                
                r_data[37132] <= r_data[37131];
                
                r_data[37133] <= r_data[37132];
                
                r_data[37134] <= r_data[37133];
                
                r_data[37135] <= r_data[37134];
                
                r_data[37136] <= r_data[37135];
                
                r_data[37137] <= r_data[37136];
                
                r_data[37138] <= r_data[37137];
                
                r_data[37139] <= r_data[37138];
                
                r_data[37140] <= r_data[37139];
                
                r_data[37141] <= r_data[37140];
                
                r_data[37142] <= r_data[37141];
                
                r_data[37143] <= r_data[37142];
                
                r_data[37144] <= r_data[37143];
                
                r_data[37145] <= r_data[37144];
                
                r_data[37146] <= r_data[37145];
                
                r_data[37147] <= r_data[37146];
                
                r_data[37148] <= r_data[37147];
                
                r_data[37149] <= r_data[37148];
                
                r_data[37150] <= r_data[37149];
                
                r_data[37151] <= r_data[37150];
                
                r_data[37152] <= r_data[37151];
                
                r_data[37153] <= r_data[37152];
                
                r_data[37154] <= r_data[37153];
                
                r_data[37155] <= r_data[37154];
                
                r_data[37156] <= r_data[37155];
                
                r_data[37157] <= r_data[37156];
                
                r_data[37158] <= r_data[37157];
                
                r_data[37159] <= r_data[37158];
                
                r_data[37160] <= r_data[37159];
                
                r_data[37161] <= r_data[37160];
                
                r_data[37162] <= r_data[37161];
                
                r_data[37163] <= r_data[37162];
                
                r_data[37164] <= r_data[37163];
                
                r_data[37165] <= r_data[37164];
                
                r_data[37166] <= r_data[37165];
                
                r_data[37167] <= r_data[37166];
                
                r_data[37168] <= r_data[37167];
                
                r_data[37169] <= r_data[37168];
                
                r_data[37170] <= r_data[37169];
                
                r_data[37171] <= r_data[37170];
                
                r_data[37172] <= r_data[37171];
                
                r_data[37173] <= r_data[37172];
                
                r_data[37174] <= r_data[37173];
                
                r_data[37175] <= r_data[37174];
                
                r_data[37176] <= r_data[37175];
                
                r_data[37177] <= r_data[37176];
                
                r_data[37178] <= r_data[37177];
                
                r_data[37179] <= r_data[37178];
                
                r_data[37180] <= r_data[37179];
                
                r_data[37181] <= r_data[37180];
                
                r_data[37182] <= r_data[37181];
                
                r_data[37183] <= r_data[37182];
                
                r_data[37184] <= r_data[37183];
                
                r_data[37185] <= r_data[37184];
                
                r_data[37186] <= r_data[37185];
                
                r_data[37187] <= r_data[37186];
                
                r_data[37188] <= r_data[37187];
                
                r_data[37189] <= r_data[37188];
                
                r_data[37190] <= r_data[37189];
                
                r_data[37191] <= r_data[37190];
                
                r_data[37192] <= r_data[37191];
                
                r_data[37193] <= r_data[37192];
                
                r_data[37194] <= r_data[37193];
                
                r_data[37195] <= r_data[37194];
                
                r_data[37196] <= r_data[37195];
                
                r_data[37197] <= r_data[37196];
                
                r_data[37198] <= r_data[37197];
                
                r_data[37199] <= r_data[37198];
                
                r_data[37200] <= r_data[37199];
                
                r_data[37201] <= r_data[37200];
                
                r_data[37202] <= r_data[37201];
                
                r_data[37203] <= r_data[37202];
                
                r_data[37204] <= r_data[37203];
                
                r_data[37205] <= r_data[37204];
                
                r_data[37206] <= r_data[37205];
                
                r_data[37207] <= r_data[37206];
                
                r_data[37208] <= r_data[37207];
                
                r_data[37209] <= r_data[37208];
                
                r_data[37210] <= r_data[37209];
                
                r_data[37211] <= r_data[37210];
                
                r_data[37212] <= r_data[37211];
                
                r_data[37213] <= r_data[37212];
                
                r_data[37214] <= r_data[37213];
                
                r_data[37215] <= r_data[37214];
                
                r_data[37216] <= r_data[37215];
                
                r_data[37217] <= r_data[37216];
                
                r_data[37218] <= r_data[37217];
                
                r_data[37219] <= r_data[37218];
                
                r_data[37220] <= r_data[37219];
                
                r_data[37221] <= r_data[37220];
                
                r_data[37222] <= r_data[37221];
                
                r_data[37223] <= r_data[37222];
                
                r_data[37224] <= r_data[37223];
                
                r_data[37225] <= r_data[37224];
                
                r_data[37226] <= r_data[37225];
                
                r_data[37227] <= r_data[37226];
                
                r_data[37228] <= r_data[37227];
                
                r_data[37229] <= r_data[37228];
                
                r_data[37230] <= r_data[37229];
                
                r_data[37231] <= r_data[37230];
                
                r_data[37232] <= r_data[37231];
                
                r_data[37233] <= r_data[37232];
                
                r_data[37234] <= r_data[37233];
                
                r_data[37235] <= r_data[37234];
                
                r_data[37236] <= r_data[37235];
                
                r_data[37237] <= r_data[37236];
                
                r_data[37238] <= r_data[37237];
                
                r_data[37239] <= r_data[37238];
                
                r_data[37240] <= r_data[37239];
                
                r_data[37241] <= r_data[37240];
                
                r_data[37242] <= r_data[37241];
                
                r_data[37243] <= r_data[37242];
                
                r_data[37244] <= r_data[37243];
                
                r_data[37245] <= r_data[37244];
                
                r_data[37246] <= r_data[37245];
                
                r_data[37247] <= r_data[37246];
                
                r_data[37248] <= r_data[37247];
                
                r_data[37249] <= r_data[37248];
                
                r_data[37250] <= r_data[37249];
                
                r_data[37251] <= r_data[37250];
                
                r_data[37252] <= r_data[37251];
                
                r_data[37253] <= r_data[37252];
                
                r_data[37254] <= r_data[37253];
                
                r_data[37255] <= r_data[37254];
                
                r_data[37256] <= r_data[37255];
                
                r_data[37257] <= r_data[37256];
                
                r_data[37258] <= r_data[37257];
                
                r_data[37259] <= r_data[37258];
                
                r_data[37260] <= r_data[37259];
                
                r_data[37261] <= r_data[37260];
                
                r_data[37262] <= r_data[37261];
                
                r_data[37263] <= r_data[37262];
                
                r_data[37264] <= r_data[37263];
                
                r_data[37265] <= r_data[37264];
                
                r_data[37266] <= r_data[37265];
                
                r_data[37267] <= r_data[37266];
                
                r_data[37268] <= r_data[37267];
                
                r_data[37269] <= r_data[37268];
                
                r_data[37270] <= r_data[37269];
                
                r_data[37271] <= r_data[37270];
                
                r_data[37272] <= r_data[37271];
                
                r_data[37273] <= r_data[37272];
                
                r_data[37274] <= r_data[37273];
                
                r_data[37275] <= r_data[37274];
                
                r_data[37276] <= r_data[37275];
                
                r_data[37277] <= r_data[37276];
                
                r_data[37278] <= r_data[37277];
                
                r_data[37279] <= r_data[37278];
                
                r_data[37280] <= r_data[37279];
                
                r_data[37281] <= r_data[37280];
                
                r_data[37282] <= r_data[37281];
                
                r_data[37283] <= r_data[37282];
                
                r_data[37284] <= r_data[37283];
                
                r_data[37285] <= r_data[37284];
                
                r_data[37286] <= r_data[37285];
                
                r_data[37287] <= r_data[37286];
                
                r_data[37288] <= r_data[37287];
                
                r_data[37289] <= r_data[37288];
                
                r_data[37290] <= r_data[37289];
                
                r_data[37291] <= r_data[37290];
                
                r_data[37292] <= r_data[37291];
                
                r_data[37293] <= r_data[37292];
                
                r_data[37294] <= r_data[37293];
                
                r_data[37295] <= r_data[37294];
                
                r_data[37296] <= r_data[37295];
                
                r_data[37297] <= r_data[37296];
                
                r_data[37298] <= r_data[37297];
                
                r_data[37299] <= r_data[37298];
                
                r_data[37300] <= r_data[37299];
                
                r_data[37301] <= r_data[37300];
                
                r_data[37302] <= r_data[37301];
                
                r_data[37303] <= r_data[37302];
                
                r_data[37304] <= r_data[37303];
                
                r_data[37305] <= r_data[37304];
                
                r_data[37306] <= r_data[37305];
                
                r_data[37307] <= r_data[37306];
                
                r_data[37308] <= r_data[37307];
                
                r_data[37309] <= r_data[37308];
                
                r_data[37310] <= r_data[37309];
                
                r_data[37311] <= r_data[37310];
                
                r_data[37312] <= r_data[37311];
                
                r_data[37313] <= r_data[37312];
                
                r_data[37314] <= r_data[37313];
                
                r_data[37315] <= r_data[37314];
                
                r_data[37316] <= r_data[37315];
                
                r_data[37317] <= r_data[37316];
                
                r_data[37318] <= r_data[37317];
                
                r_data[37319] <= r_data[37318];
                
                r_data[37320] <= r_data[37319];
                
                r_data[37321] <= r_data[37320];
                
                r_data[37322] <= r_data[37321];
                
                r_data[37323] <= r_data[37322];
                
                r_data[37324] <= r_data[37323];
                
                r_data[37325] <= r_data[37324];
                
                r_data[37326] <= r_data[37325];
                
                r_data[37327] <= r_data[37326];
                
                r_data[37328] <= r_data[37327];
                
                r_data[37329] <= r_data[37328];
                
                r_data[37330] <= r_data[37329];
                
                r_data[37331] <= r_data[37330];
                
                r_data[37332] <= r_data[37331];
                
                r_data[37333] <= r_data[37332];
                
                r_data[37334] <= r_data[37333];
                
                r_data[37335] <= r_data[37334];
                
                r_data[37336] <= r_data[37335];
                
                r_data[37337] <= r_data[37336];
                
                r_data[37338] <= r_data[37337];
                
                r_data[37339] <= r_data[37338];
                
                r_data[37340] <= r_data[37339];
                
                r_data[37341] <= r_data[37340];
                
                r_data[37342] <= r_data[37341];
                
                r_data[37343] <= r_data[37342];
                
                r_data[37344] <= r_data[37343];
                
                r_data[37345] <= r_data[37344];
                
                r_data[37346] <= r_data[37345];
                
                r_data[37347] <= r_data[37346];
                
                r_data[37348] <= r_data[37347];
                
                r_data[37349] <= r_data[37348];
                
                r_data[37350] <= r_data[37349];
                
                r_data[37351] <= r_data[37350];
                
                r_data[37352] <= r_data[37351];
                
                r_data[37353] <= r_data[37352];
                
                r_data[37354] <= r_data[37353];
                
                r_data[37355] <= r_data[37354];
                
                r_data[37356] <= r_data[37355];
                
                r_data[37357] <= r_data[37356];
                
                r_data[37358] <= r_data[37357];
                
                r_data[37359] <= r_data[37358];
                
                r_data[37360] <= r_data[37359];
                
                r_data[37361] <= r_data[37360];
                
                r_data[37362] <= r_data[37361];
                
                r_data[37363] <= r_data[37362];
                
                r_data[37364] <= r_data[37363];
                
                r_data[37365] <= r_data[37364];
                
                r_data[37366] <= r_data[37365];
                
                r_data[37367] <= r_data[37366];
                
                r_data[37368] <= r_data[37367];
                
                r_data[37369] <= r_data[37368];
                
                r_data[37370] <= r_data[37369];
                
                r_data[37371] <= r_data[37370];
                
                r_data[37372] <= r_data[37371];
                
                r_data[37373] <= r_data[37372];
                
                r_data[37374] <= r_data[37373];
                
                r_data[37375] <= r_data[37374];
                
                r_data[37376] <= r_data[37375];
                
                r_data[37377] <= r_data[37376];
                
                r_data[37378] <= r_data[37377];
                
                r_data[37379] <= r_data[37378];
                
                r_data[37380] <= r_data[37379];
                
                r_data[37381] <= r_data[37380];
                
                r_data[37382] <= r_data[37381];
                
                r_data[37383] <= r_data[37382];
                
                r_data[37384] <= r_data[37383];
                
                r_data[37385] <= r_data[37384];
                
                r_data[37386] <= r_data[37385];
                
                r_data[37387] <= r_data[37386];
                
                r_data[37388] <= r_data[37387];
                
                r_data[37389] <= r_data[37388];
                
                r_data[37390] <= r_data[37389];
                
                r_data[37391] <= r_data[37390];
                
                r_data[37392] <= r_data[37391];
                
                r_data[37393] <= r_data[37392];
                
                r_data[37394] <= r_data[37393];
                
                r_data[37395] <= r_data[37394];
                
                r_data[37396] <= r_data[37395];
                
                r_data[37397] <= r_data[37396];
                
                r_data[37398] <= r_data[37397];
                
                r_data[37399] <= r_data[37398];
                
                r_data[37400] <= r_data[37399];
                
                r_data[37401] <= r_data[37400];
                
                r_data[37402] <= r_data[37401];
                
                r_data[37403] <= r_data[37402];
                
                r_data[37404] <= r_data[37403];
                
                r_data[37405] <= r_data[37404];
                
                r_data[37406] <= r_data[37405];
                
                r_data[37407] <= r_data[37406];
                
                r_data[37408] <= r_data[37407];
                
                r_data[37409] <= r_data[37408];
                
                r_data[37410] <= r_data[37409];
                
                r_data[37411] <= r_data[37410];
                
                r_data[37412] <= r_data[37411];
                
                r_data[37413] <= r_data[37412];
                
                r_data[37414] <= r_data[37413];
                
                r_data[37415] <= r_data[37414];
                
                r_data[37416] <= r_data[37415];
                
                r_data[37417] <= r_data[37416];
                
                r_data[37418] <= r_data[37417];
                
                r_data[37419] <= r_data[37418];
                
                r_data[37420] <= r_data[37419];
                
                r_data[37421] <= r_data[37420];
                
                r_data[37422] <= r_data[37421];
                
                r_data[37423] <= r_data[37422];
                
                r_data[37424] <= r_data[37423];
                
                r_data[37425] <= r_data[37424];
                
                r_data[37426] <= r_data[37425];
                
                r_data[37427] <= r_data[37426];
                
                r_data[37428] <= r_data[37427];
                
                r_data[37429] <= r_data[37428];
                
                r_data[37430] <= r_data[37429];
                
                r_data[37431] <= r_data[37430];
                
                r_data[37432] <= r_data[37431];
                
                r_data[37433] <= r_data[37432];
                
                r_data[37434] <= r_data[37433];
                
                r_data[37435] <= r_data[37434];
                
                r_data[37436] <= r_data[37435];
                
                r_data[37437] <= r_data[37436];
                
                r_data[37438] <= r_data[37437];
                
                r_data[37439] <= r_data[37438];
                
                r_data[37440] <= r_data[37439];
                
                r_data[37441] <= r_data[37440];
                
                r_data[37442] <= r_data[37441];
                
                r_data[37443] <= r_data[37442];
                
                r_data[37444] <= r_data[37443];
                
                r_data[37445] <= r_data[37444];
                
                r_data[37446] <= r_data[37445];
                
                r_data[37447] <= r_data[37446];
                
                r_data[37448] <= r_data[37447];
                
                r_data[37449] <= r_data[37448];
                
                r_data[37450] <= r_data[37449];
                
                r_data[37451] <= r_data[37450];
                
                r_data[37452] <= r_data[37451];
                
                r_data[37453] <= r_data[37452];
                
                r_data[37454] <= r_data[37453];
                
                r_data[37455] <= r_data[37454];
                
                r_data[37456] <= r_data[37455];
                
                r_data[37457] <= r_data[37456];
                
                r_data[37458] <= r_data[37457];
                
                r_data[37459] <= r_data[37458];
                
                r_data[37460] <= r_data[37459];
                
                r_data[37461] <= r_data[37460];
                
                r_data[37462] <= r_data[37461];
                
                r_data[37463] <= r_data[37462];
                
                r_data[37464] <= r_data[37463];
                
                r_data[37465] <= r_data[37464];
                
                r_data[37466] <= r_data[37465];
                
                r_data[37467] <= r_data[37466];
                
                r_data[37468] <= r_data[37467];
                
                r_data[37469] <= r_data[37468];
                
                r_data[37470] <= r_data[37469];
                
                r_data[37471] <= r_data[37470];
                
                r_data[37472] <= r_data[37471];
                
                r_data[37473] <= r_data[37472];
                
                r_data[37474] <= r_data[37473];
                
                r_data[37475] <= r_data[37474];
                
                r_data[37476] <= r_data[37475];
                
                r_data[37477] <= r_data[37476];
                
                r_data[37478] <= r_data[37477];
                
                r_data[37479] <= r_data[37478];
                
                r_data[37480] <= r_data[37479];
                
                r_data[37481] <= r_data[37480];
                
                r_data[37482] <= r_data[37481];
                
                r_data[37483] <= r_data[37482];
                
                r_data[37484] <= r_data[37483];
                
                r_data[37485] <= r_data[37484];
                
                r_data[37486] <= r_data[37485];
                
                r_data[37487] <= r_data[37486];
                
                r_data[37488] <= r_data[37487];
                
                r_data[37489] <= r_data[37488];
                
                r_data[37490] <= r_data[37489];
                
                r_data[37491] <= r_data[37490];
                
                r_data[37492] <= r_data[37491];
                
                r_data[37493] <= r_data[37492];
                
                r_data[37494] <= r_data[37493];
                
                r_data[37495] <= r_data[37494];
                
                r_data[37496] <= r_data[37495];
                
                r_data[37497] <= r_data[37496];
                
                r_data[37498] <= r_data[37497];
                
                r_data[37499] <= r_data[37498];
                
                r_data[37500] <= r_data[37499];
                
                r_data[37501] <= r_data[37500];
                
                r_data[37502] <= r_data[37501];
                
                r_data[37503] <= r_data[37502];
                
                r_data[37504] <= r_data[37503];
                
                r_data[37505] <= r_data[37504];
                
                r_data[37506] <= r_data[37505];
                
                r_data[37507] <= r_data[37506];
                
                r_data[37508] <= r_data[37507];
                
                r_data[37509] <= r_data[37508];
                
                r_data[37510] <= r_data[37509];
                
                r_data[37511] <= r_data[37510];
                
                r_data[37512] <= r_data[37511];
                
                r_data[37513] <= r_data[37512];
                
                r_data[37514] <= r_data[37513];
                
                r_data[37515] <= r_data[37514];
                
                r_data[37516] <= r_data[37515];
                
                r_data[37517] <= r_data[37516];
                
                r_data[37518] <= r_data[37517];
                
                r_data[37519] <= r_data[37518];
                
                r_data[37520] <= r_data[37519];
                
                r_data[37521] <= r_data[37520];
                
                r_data[37522] <= r_data[37521];
                
                r_data[37523] <= r_data[37522];
                
                r_data[37524] <= r_data[37523];
                
                r_data[37525] <= r_data[37524];
                
                r_data[37526] <= r_data[37525];
                
                r_data[37527] <= r_data[37526];
                
                r_data[37528] <= r_data[37527];
                
                r_data[37529] <= r_data[37528];
                
                r_data[37530] <= r_data[37529];
                
                r_data[37531] <= r_data[37530];
                
                r_data[37532] <= r_data[37531];
                
                r_data[37533] <= r_data[37532];
                
                r_data[37534] <= r_data[37533];
                
                r_data[37535] <= r_data[37534];
                
                r_data[37536] <= r_data[37535];
                
                r_data[37537] <= r_data[37536];
                
                r_data[37538] <= r_data[37537];
                
                r_data[37539] <= r_data[37538];
                
                r_data[37540] <= r_data[37539];
                
                r_data[37541] <= r_data[37540];
                
                r_data[37542] <= r_data[37541];
                
                r_data[37543] <= r_data[37542];
                
                r_data[37544] <= r_data[37543];
                
                r_data[37545] <= r_data[37544];
                
                r_data[37546] <= r_data[37545];
                
                r_data[37547] <= r_data[37546];
                
                r_data[37548] <= r_data[37547];
                
                r_data[37549] <= r_data[37548];
                
                r_data[37550] <= r_data[37549];
                
                r_data[37551] <= r_data[37550];
                
                r_data[37552] <= r_data[37551];
                
                r_data[37553] <= r_data[37552];
                
                r_data[37554] <= r_data[37553];
                
                r_data[37555] <= r_data[37554];
                
                r_data[37556] <= r_data[37555];
                
                r_data[37557] <= r_data[37556];
                
                r_data[37558] <= r_data[37557];
                
                r_data[37559] <= r_data[37558];
                
                r_data[37560] <= r_data[37559];
                
                r_data[37561] <= r_data[37560];
                
                r_data[37562] <= r_data[37561];
                
                r_data[37563] <= r_data[37562];
                
                r_data[37564] <= r_data[37563];
                
                r_data[37565] <= r_data[37564];
                
                r_data[37566] <= r_data[37565];
                
                r_data[37567] <= r_data[37566];
                
                r_data[37568] <= r_data[37567];
                
                r_data[37569] <= r_data[37568];
                
                r_data[37570] <= r_data[37569];
                
                r_data[37571] <= r_data[37570];
                
                r_data[37572] <= r_data[37571];
                
                r_data[37573] <= r_data[37572];
                
                r_data[37574] <= r_data[37573];
                
                r_data[37575] <= r_data[37574];
                
                r_data[37576] <= r_data[37575];
                
                r_data[37577] <= r_data[37576];
                
                r_data[37578] <= r_data[37577];
                
                r_data[37579] <= r_data[37578];
                
                r_data[37580] <= r_data[37579];
                
                r_data[37581] <= r_data[37580];
                
                r_data[37582] <= r_data[37581];
                
                r_data[37583] <= r_data[37582];
                
                r_data[37584] <= r_data[37583];
                
                r_data[37585] <= r_data[37584];
                
                r_data[37586] <= r_data[37585];
                
                r_data[37587] <= r_data[37586];
                
                r_data[37588] <= r_data[37587];
                
                r_data[37589] <= r_data[37588];
                
                r_data[37590] <= r_data[37589];
                
                r_data[37591] <= r_data[37590];
                
                r_data[37592] <= r_data[37591];
                
                r_data[37593] <= r_data[37592];
                
                r_data[37594] <= r_data[37593];
                
                r_data[37595] <= r_data[37594];
                
                r_data[37596] <= r_data[37595];
                
                r_data[37597] <= r_data[37596];
                
                r_data[37598] <= r_data[37597];
                
                r_data[37599] <= r_data[37598];
                
                r_data[37600] <= r_data[37599];
                
                r_data[37601] <= r_data[37600];
                
                r_data[37602] <= r_data[37601];
                
                r_data[37603] <= r_data[37602];
                
                r_data[37604] <= r_data[37603];
                
                r_data[37605] <= r_data[37604];
                
                r_data[37606] <= r_data[37605];
                
                r_data[37607] <= r_data[37606];
                
                r_data[37608] <= r_data[37607];
                
                r_data[37609] <= r_data[37608];
                
                r_data[37610] <= r_data[37609];
                
                r_data[37611] <= r_data[37610];
                
                r_data[37612] <= r_data[37611];
                
                r_data[37613] <= r_data[37612];
                
                r_data[37614] <= r_data[37613];
                
                r_data[37615] <= r_data[37614];
                
                r_data[37616] <= r_data[37615];
                
                r_data[37617] <= r_data[37616];
                
                r_data[37618] <= r_data[37617];
                
                r_data[37619] <= r_data[37618];
                
                r_data[37620] <= r_data[37619];
                
                r_data[37621] <= r_data[37620];
                
                r_data[37622] <= r_data[37621];
                
                r_data[37623] <= r_data[37622];
                
                r_data[37624] <= r_data[37623];
                
                r_data[37625] <= r_data[37624];
                
                r_data[37626] <= r_data[37625];
                
                r_data[37627] <= r_data[37626];
                
                r_data[37628] <= r_data[37627];
                
                r_data[37629] <= r_data[37628];
                
                r_data[37630] <= r_data[37629];
                
                r_data[37631] <= r_data[37630];
                
                r_data[37632] <= r_data[37631];
                
                r_data[37633] <= r_data[37632];
                
                r_data[37634] <= r_data[37633];
                
                r_data[37635] <= r_data[37634];
                
                r_data[37636] <= r_data[37635];
                
                r_data[37637] <= r_data[37636];
                
                r_data[37638] <= r_data[37637];
                
                r_data[37639] <= r_data[37638];
                
                r_data[37640] <= r_data[37639];
                
                r_data[37641] <= r_data[37640];
                
                r_data[37642] <= r_data[37641];
                
                r_data[37643] <= r_data[37642];
                
                r_data[37644] <= r_data[37643];
                
                r_data[37645] <= r_data[37644];
                
                r_data[37646] <= r_data[37645];
                
                r_data[37647] <= r_data[37646];
                
                r_data[37648] <= r_data[37647];
                
                r_data[37649] <= r_data[37648];
                
                r_data[37650] <= r_data[37649];
                
                r_data[37651] <= r_data[37650];
                
                r_data[37652] <= r_data[37651];
                
                r_data[37653] <= r_data[37652];
                
                r_data[37654] <= r_data[37653];
                
                r_data[37655] <= r_data[37654];
                
                r_data[37656] <= r_data[37655];
                
                r_data[37657] <= r_data[37656];
                
                r_data[37658] <= r_data[37657];
                
                r_data[37659] <= r_data[37658];
                
                r_data[37660] <= r_data[37659];
                
                r_data[37661] <= r_data[37660];
                
                r_data[37662] <= r_data[37661];
                
                r_data[37663] <= r_data[37662];
                
                r_data[37664] <= r_data[37663];
                
                r_data[37665] <= r_data[37664];
                
                r_data[37666] <= r_data[37665];
                
                r_data[37667] <= r_data[37666];
                
                r_data[37668] <= r_data[37667];
                
                r_data[37669] <= r_data[37668];
                
                r_data[37670] <= r_data[37669];
                
                r_data[37671] <= r_data[37670];
                
                r_data[37672] <= r_data[37671];
                
                r_data[37673] <= r_data[37672];
                
                r_data[37674] <= r_data[37673];
                
                r_data[37675] <= r_data[37674];
                
                r_data[37676] <= r_data[37675];
                
                r_data[37677] <= r_data[37676];
                
                r_data[37678] <= r_data[37677];
                
                r_data[37679] <= r_data[37678];
                
                r_data[37680] <= r_data[37679];
                
                r_data[37681] <= r_data[37680];
                
                r_data[37682] <= r_data[37681];
                
                r_data[37683] <= r_data[37682];
                
                r_data[37684] <= r_data[37683];
                
                r_data[37685] <= r_data[37684];
                
                r_data[37686] <= r_data[37685];
                
                r_data[37687] <= r_data[37686];
                
                r_data[37688] <= r_data[37687];
                
                r_data[37689] <= r_data[37688];
                
                r_data[37690] <= r_data[37689];
                
                r_data[37691] <= r_data[37690];
                
                r_data[37692] <= r_data[37691];
                
                r_data[37693] <= r_data[37692];
                
                r_data[37694] <= r_data[37693];
                
                r_data[37695] <= r_data[37694];
                
                r_data[37696] <= r_data[37695];
                
                r_data[37697] <= r_data[37696];
                
                r_data[37698] <= r_data[37697];
                
                r_data[37699] <= r_data[37698];
                
                r_data[37700] <= r_data[37699];
                
                r_data[37701] <= r_data[37700];
                
                r_data[37702] <= r_data[37701];
                
                r_data[37703] <= r_data[37702];
                
                r_data[37704] <= r_data[37703];
                
                r_data[37705] <= r_data[37704];
                
                r_data[37706] <= r_data[37705];
                
                r_data[37707] <= r_data[37706];
                
                r_data[37708] <= r_data[37707];
                
                r_data[37709] <= r_data[37708];
                
                r_data[37710] <= r_data[37709];
                
                r_data[37711] <= r_data[37710];
                
                r_data[37712] <= r_data[37711];
                
                r_data[37713] <= r_data[37712];
                
                r_data[37714] <= r_data[37713];
                
                r_data[37715] <= r_data[37714];
                
                r_data[37716] <= r_data[37715];
                
                r_data[37717] <= r_data[37716];
                
                r_data[37718] <= r_data[37717];
                
                r_data[37719] <= r_data[37718];
                
                r_data[37720] <= r_data[37719];
                
                r_data[37721] <= r_data[37720];
                
                r_data[37722] <= r_data[37721];
                
                r_data[37723] <= r_data[37722];
                
                r_data[37724] <= r_data[37723];
                
                r_data[37725] <= r_data[37724];
                
                r_data[37726] <= r_data[37725];
                
                r_data[37727] <= r_data[37726];
                
                r_data[37728] <= r_data[37727];
                
                r_data[37729] <= r_data[37728];
                
                r_data[37730] <= r_data[37729];
                
                r_data[37731] <= r_data[37730];
                
                r_data[37732] <= r_data[37731];
                
                r_data[37733] <= r_data[37732];
                
                r_data[37734] <= r_data[37733];
                
                r_data[37735] <= r_data[37734];
                
                r_data[37736] <= r_data[37735];
                
                r_data[37737] <= r_data[37736];
                
                r_data[37738] <= r_data[37737];
                
                r_data[37739] <= r_data[37738];
                
                r_data[37740] <= r_data[37739];
                
                r_data[37741] <= r_data[37740];
                
                r_data[37742] <= r_data[37741];
                
                r_data[37743] <= r_data[37742];
                
                r_data[37744] <= r_data[37743];
                
                r_data[37745] <= r_data[37744];
                
                r_data[37746] <= r_data[37745];
                
                r_data[37747] <= r_data[37746];
                
                r_data[37748] <= r_data[37747];
                
                r_data[37749] <= r_data[37748];
                
                r_data[37750] <= r_data[37749];
                
                r_data[37751] <= r_data[37750];
                
                r_data[37752] <= r_data[37751];
                
                r_data[37753] <= r_data[37752];
                
                r_data[37754] <= r_data[37753];
                
                r_data[37755] <= r_data[37754];
                
                r_data[37756] <= r_data[37755];
                
                r_data[37757] <= r_data[37756];
                
                r_data[37758] <= r_data[37757];
                
                r_data[37759] <= r_data[37758];
                
                r_data[37760] <= r_data[37759];
                
                r_data[37761] <= r_data[37760];
                
                r_data[37762] <= r_data[37761];
                
                r_data[37763] <= r_data[37762];
                
                r_data[37764] <= r_data[37763];
                
                r_data[37765] <= r_data[37764];
                
                r_data[37766] <= r_data[37765];
                
                r_data[37767] <= r_data[37766];
                
                r_data[37768] <= r_data[37767];
                
                r_data[37769] <= r_data[37768];
                
                r_data[37770] <= r_data[37769];
                
                r_data[37771] <= r_data[37770];
                
                r_data[37772] <= r_data[37771];
                
                r_data[37773] <= r_data[37772];
                
                r_data[37774] <= r_data[37773];
                
                r_data[37775] <= r_data[37774];
                
                r_data[37776] <= r_data[37775];
                
                r_data[37777] <= r_data[37776];
                
                r_data[37778] <= r_data[37777];
                
                r_data[37779] <= r_data[37778];
                
                r_data[37780] <= r_data[37779];
                
                r_data[37781] <= r_data[37780];
                
                r_data[37782] <= r_data[37781];
                
                r_data[37783] <= r_data[37782];
                
                r_data[37784] <= r_data[37783];
                
                r_data[37785] <= r_data[37784];
                
                r_data[37786] <= r_data[37785];
                
                r_data[37787] <= r_data[37786];
                
                r_data[37788] <= r_data[37787];
                
                r_data[37789] <= r_data[37788];
                
                r_data[37790] <= r_data[37789];
                
                r_data[37791] <= r_data[37790];
                
                r_data[37792] <= r_data[37791];
                
                r_data[37793] <= r_data[37792];
                
                r_data[37794] <= r_data[37793];
                
                r_data[37795] <= r_data[37794];
                
                r_data[37796] <= r_data[37795];
                
                r_data[37797] <= r_data[37796];
                
                r_data[37798] <= r_data[37797];
                
                r_data[37799] <= r_data[37798];
                
                r_data[37800] <= r_data[37799];
                
                r_data[37801] <= r_data[37800];
                
                r_data[37802] <= r_data[37801];
                
                r_data[37803] <= r_data[37802];
                
                r_data[37804] <= r_data[37803];
                
                r_data[37805] <= r_data[37804];
                
                r_data[37806] <= r_data[37805];
                
                r_data[37807] <= r_data[37806];
                
                r_data[37808] <= r_data[37807];
                
                r_data[37809] <= r_data[37808];
                
                r_data[37810] <= r_data[37809];
                
                r_data[37811] <= r_data[37810];
                
                r_data[37812] <= r_data[37811];
                
                r_data[37813] <= r_data[37812];
                
                r_data[37814] <= r_data[37813];
                
                r_data[37815] <= r_data[37814];
                
                r_data[37816] <= r_data[37815];
                
                r_data[37817] <= r_data[37816];
                
                r_data[37818] <= r_data[37817];
                
                r_data[37819] <= r_data[37818];
                
                r_data[37820] <= r_data[37819];
                
                r_data[37821] <= r_data[37820];
                
                r_data[37822] <= r_data[37821];
                
                r_data[37823] <= r_data[37822];
                
                r_data[37824] <= r_data[37823];
                
                r_data[37825] <= r_data[37824];
                
                r_data[37826] <= r_data[37825];
                
                r_data[37827] <= r_data[37826];
                
                r_data[37828] <= r_data[37827];
                
                r_data[37829] <= r_data[37828];
                
                r_data[37830] <= r_data[37829];
                
                r_data[37831] <= r_data[37830];
                
                r_data[37832] <= r_data[37831];
                
                r_data[37833] <= r_data[37832];
                
                r_data[37834] <= r_data[37833];
                
                r_data[37835] <= r_data[37834];
                
                r_data[37836] <= r_data[37835];
                
                r_data[37837] <= r_data[37836];
                
                r_data[37838] <= r_data[37837];
                
                r_data[37839] <= r_data[37838];
                
                r_data[37840] <= r_data[37839];
                
                r_data[37841] <= r_data[37840];
                
                r_data[37842] <= r_data[37841];
                
                r_data[37843] <= r_data[37842];
                
                r_data[37844] <= r_data[37843];
                
                r_data[37845] <= r_data[37844];
                
                r_data[37846] <= r_data[37845];
                
                r_data[37847] <= r_data[37846];
                
                r_data[37848] <= r_data[37847];
                
                r_data[37849] <= r_data[37848];
                
                r_data[37850] <= r_data[37849];
                
                r_data[37851] <= r_data[37850];
                
                r_data[37852] <= r_data[37851];
                
                r_data[37853] <= r_data[37852];
                
                r_data[37854] <= r_data[37853];
                
                r_data[37855] <= r_data[37854];
                
                r_data[37856] <= r_data[37855];
                
                r_data[37857] <= r_data[37856];
                
                r_data[37858] <= r_data[37857];
                
                r_data[37859] <= r_data[37858];
                
                r_data[37860] <= r_data[37859];
                
                r_data[37861] <= r_data[37860];
                
                r_data[37862] <= r_data[37861];
                
                r_data[37863] <= r_data[37862];
                
                r_data[37864] <= r_data[37863];
                
                r_data[37865] <= r_data[37864];
                
                r_data[37866] <= r_data[37865];
                
                r_data[37867] <= r_data[37866];
                
                r_data[37868] <= r_data[37867];
                
                r_data[37869] <= r_data[37868];
                
                r_data[37870] <= r_data[37869];
                
                r_data[37871] <= r_data[37870];
                
                r_data[37872] <= r_data[37871];
                
                r_data[37873] <= r_data[37872];
                
                r_data[37874] <= r_data[37873];
                
                r_data[37875] <= r_data[37874];
                
                r_data[37876] <= r_data[37875];
                
                r_data[37877] <= r_data[37876];
                
                r_data[37878] <= r_data[37877];
                
                r_data[37879] <= r_data[37878];
                
                r_data[37880] <= r_data[37879];
                
                r_data[37881] <= r_data[37880];
                
                r_data[37882] <= r_data[37881];
                
                r_data[37883] <= r_data[37882];
                
                r_data[37884] <= r_data[37883];
                
                r_data[37885] <= r_data[37884];
                
                r_data[37886] <= r_data[37885];
                
                r_data[37887] <= r_data[37886];
                
                r_data[37888] <= r_data[37887];
                
                r_data[37889] <= r_data[37888];
                
                r_data[37890] <= r_data[37889];
                
                r_data[37891] <= r_data[37890];
                
                r_data[37892] <= r_data[37891];
                
                r_data[37893] <= r_data[37892];
                
                r_data[37894] <= r_data[37893];
                
                r_data[37895] <= r_data[37894];
                
                r_data[37896] <= r_data[37895];
                
                r_data[37897] <= r_data[37896];
                
                r_data[37898] <= r_data[37897];
                
                r_data[37899] <= r_data[37898];
                
                r_data[37900] <= r_data[37899];
                
                r_data[37901] <= r_data[37900];
                
                r_data[37902] <= r_data[37901];
                
                r_data[37903] <= r_data[37902];
                
                r_data[37904] <= r_data[37903];
                
                r_data[37905] <= r_data[37904];
                
                r_data[37906] <= r_data[37905];
                
                r_data[37907] <= r_data[37906];
                
                r_data[37908] <= r_data[37907];
                
                r_data[37909] <= r_data[37908];
                
                r_data[37910] <= r_data[37909];
                
                r_data[37911] <= r_data[37910];
                
                r_data[37912] <= r_data[37911];
                
                r_data[37913] <= r_data[37912];
                
                r_data[37914] <= r_data[37913];
                
                r_data[37915] <= r_data[37914];
                
                r_data[37916] <= r_data[37915];
                
                r_data[37917] <= r_data[37916];
                
                r_data[37918] <= r_data[37917];
                
                r_data[37919] <= r_data[37918];
                
                r_data[37920] <= r_data[37919];
                
                r_data[37921] <= r_data[37920];
                
                r_data[37922] <= r_data[37921];
                
                r_data[37923] <= r_data[37922];
                
                r_data[37924] <= r_data[37923];
                
                r_data[37925] <= r_data[37924];
                
                r_data[37926] <= r_data[37925];
                
                r_data[37927] <= r_data[37926];
                
                r_data[37928] <= r_data[37927];
                
                r_data[37929] <= r_data[37928];
                
                r_data[37930] <= r_data[37929];
                
                r_data[37931] <= r_data[37930];
                
                r_data[37932] <= r_data[37931];
                
                r_data[37933] <= r_data[37932];
                
                r_data[37934] <= r_data[37933];
                
                r_data[37935] <= r_data[37934];
                
                r_data[37936] <= r_data[37935];
                
                r_data[37937] <= r_data[37936];
                
                r_data[37938] <= r_data[37937];
                
                r_data[37939] <= r_data[37938];
                
                r_data[37940] <= r_data[37939];
                
                r_data[37941] <= r_data[37940];
                
                r_data[37942] <= r_data[37941];
                
                r_data[37943] <= r_data[37942];
                
                r_data[37944] <= r_data[37943];
                
                r_data[37945] <= r_data[37944];
                
                r_data[37946] <= r_data[37945];
                
                r_data[37947] <= r_data[37946];
                
                r_data[37948] <= r_data[37947];
                
                r_data[37949] <= r_data[37948];
                
                r_data[37950] <= r_data[37949];
                
                r_data[37951] <= r_data[37950];
                
                r_data[37952] <= r_data[37951];
                
                r_data[37953] <= r_data[37952];
                
                r_data[37954] <= r_data[37953];
                
                r_data[37955] <= r_data[37954];
                
                r_data[37956] <= r_data[37955];
                
                r_data[37957] <= r_data[37956];
                
                r_data[37958] <= r_data[37957];
                
                r_data[37959] <= r_data[37958];
                
                r_data[37960] <= r_data[37959];
                
                r_data[37961] <= r_data[37960];
                
                r_data[37962] <= r_data[37961];
                
                r_data[37963] <= r_data[37962];
                
                r_data[37964] <= r_data[37963];
                
                r_data[37965] <= r_data[37964];
                
                r_data[37966] <= r_data[37965];
                
                r_data[37967] <= r_data[37966];
                
                r_data[37968] <= r_data[37967];
                
                r_data[37969] <= r_data[37968];
                
                r_data[37970] <= r_data[37969];
                
                r_data[37971] <= r_data[37970];
                
                r_data[37972] <= r_data[37971];
                
                r_data[37973] <= r_data[37972];
                
                r_data[37974] <= r_data[37973];
                
                r_data[37975] <= r_data[37974];
                
                r_data[37976] <= r_data[37975];
                
                r_data[37977] <= r_data[37976];
                
                r_data[37978] <= r_data[37977];
                
                r_data[37979] <= r_data[37978];
                
                r_data[37980] <= r_data[37979];
                
                r_data[37981] <= r_data[37980];
                
                r_data[37982] <= r_data[37981];
                
                r_data[37983] <= r_data[37982];
                
                r_data[37984] <= r_data[37983];
                
                r_data[37985] <= r_data[37984];
                
                r_data[37986] <= r_data[37985];
                
                r_data[37987] <= r_data[37986];
                
                r_data[37988] <= r_data[37987];
                
                r_data[37989] <= r_data[37988];
                
                r_data[37990] <= r_data[37989];
                
                r_data[37991] <= r_data[37990];
                
                r_data[37992] <= r_data[37991];
                
                r_data[37993] <= r_data[37992];
                
                r_data[37994] <= r_data[37993];
                
                r_data[37995] <= r_data[37994];
                
                r_data[37996] <= r_data[37995];
                
                r_data[37997] <= r_data[37996];
                
                r_data[37998] <= r_data[37997];
                
                r_data[37999] <= r_data[37998];
                
                r_data[38000] <= r_data[37999];
                
                r_data[38001] <= r_data[38000];
                
                r_data[38002] <= r_data[38001];
                
                r_data[38003] <= r_data[38002];
                
                r_data[38004] <= r_data[38003];
                
                r_data[38005] <= r_data[38004];
                
                r_data[38006] <= r_data[38005];
                
                r_data[38007] <= r_data[38006];
                
                r_data[38008] <= r_data[38007];
                
                r_data[38009] <= r_data[38008];
                
                r_data[38010] <= r_data[38009];
                
                r_data[38011] <= r_data[38010];
                
                r_data[38012] <= r_data[38011];
                
                r_data[38013] <= r_data[38012];
                
                r_data[38014] <= r_data[38013];
                
                r_data[38015] <= r_data[38014];
                
                r_data[38016] <= r_data[38015];
                
                r_data[38017] <= r_data[38016];
                
                r_data[38018] <= r_data[38017];
                
                r_data[38019] <= r_data[38018];
                
                r_data[38020] <= r_data[38019];
                
                r_data[38021] <= r_data[38020];
                
                r_data[38022] <= r_data[38021];
                
                r_data[38023] <= r_data[38022];
                
                r_data[38024] <= r_data[38023];
                
                r_data[38025] <= r_data[38024];
                
                r_data[38026] <= r_data[38025];
                
                r_data[38027] <= r_data[38026];
                
                r_data[38028] <= r_data[38027];
                
                r_data[38029] <= r_data[38028];
                
                r_data[38030] <= r_data[38029];
                
                r_data[38031] <= r_data[38030];
                
                r_data[38032] <= r_data[38031];
                
                r_data[38033] <= r_data[38032];
                
                r_data[38034] <= r_data[38033];
                
                r_data[38035] <= r_data[38034];
                
                r_data[38036] <= r_data[38035];
                
                r_data[38037] <= r_data[38036];
                
                r_data[38038] <= r_data[38037];
                
                r_data[38039] <= r_data[38038];
                
                r_data[38040] <= r_data[38039];
                
                r_data[38041] <= r_data[38040];
                
                r_data[38042] <= r_data[38041];
                
                r_data[38043] <= r_data[38042];
                
                r_data[38044] <= r_data[38043];
                
                r_data[38045] <= r_data[38044];
                
                r_data[38046] <= r_data[38045];
                
                r_data[38047] <= r_data[38046];
                
                r_data[38048] <= r_data[38047];
                
                r_data[38049] <= r_data[38048];
                
                r_data[38050] <= r_data[38049];
                
                r_data[38051] <= r_data[38050];
                
                r_data[38052] <= r_data[38051];
                
                r_data[38053] <= r_data[38052];
                
                r_data[38054] <= r_data[38053];
                
                r_data[38055] <= r_data[38054];
                
                r_data[38056] <= r_data[38055];
                
                r_data[38057] <= r_data[38056];
                
                r_data[38058] <= r_data[38057];
                
                r_data[38059] <= r_data[38058];
                
                r_data[38060] <= r_data[38059];
                
                r_data[38061] <= r_data[38060];
                
                r_data[38062] <= r_data[38061];
                
                r_data[38063] <= r_data[38062];
                
                r_data[38064] <= r_data[38063];
                
                r_data[38065] <= r_data[38064];
                
                r_data[38066] <= r_data[38065];
                
                r_data[38067] <= r_data[38066];
                
                r_data[38068] <= r_data[38067];
                
                r_data[38069] <= r_data[38068];
                
                r_data[38070] <= r_data[38069];
                
                r_data[38071] <= r_data[38070];
                
                r_data[38072] <= r_data[38071];
                
                r_data[38073] <= r_data[38072];
                
                r_data[38074] <= r_data[38073];
                
                r_data[38075] <= r_data[38074];
                
                r_data[38076] <= r_data[38075];
                
                r_data[38077] <= r_data[38076];
                
                r_data[38078] <= r_data[38077];
                
                r_data[38079] <= r_data[38078];
                
                r_data[38080] <= r_data[38079];
                
                r_data[38081] <= r_data[38080];
                
                r_data[38082] <= r_data[38081];
                
                r_data[38083] <= r_data[38082];
                
                r_data[38084] <= r_data[38083];
                
                r_data[38085] <= r_data[38084];
                
                r_data[38086] <= r_data[38085];
                
                r_data[38087] <= r_data[38086];
                
                r_data[38088] <= r_data[38087];
                
                r_data[38089] <= r_data[38088];
                
                r_data[38090] <= r_data[38089];
                
                r_data[38091] <= r_data[38090];
                
                r_data[38092] <= r_data[38091];
                
                r_data[38093] <= r_data[38092];
                
                r_data[38094] <= r_data[38093];
                
                r_data[38095] <= r_data[38094];
                
                r_data[38096] <= r_data[38095];
                
                r_data[38097] <= r_data[38096];
                
                r_data[38098] <= r_data[38097];
                
                r_data[38099] <= r_data[38098];
                
                r_data[38100] <= r_data[38099];
                
                r_data[38101] <= r_data[38100];
                
                r_data[38102] <= r_data[38101];
                
                r_data[38103] <= r_data[38102];
                
                r_data[38104] <= r_data[38103];
                
                r_data[38105] <= r_data[38104];
                
                r_data[38106] <= r_data[38105];
                
                r_data[38107] <= r_data[38106];
                
                r_data[38108] <= r_data[38107];
                
                r_data[38109] <= r_data[38108];
                
                r_data[38110] <= r_data[38109];
                
                r_data[38111] <= r_data[38110];
                
                r_data[38112] <= r_data[38111];
                
                r_data[38113] <= r_data[38112];
                
                r_data[38114] <= r_data[38113];
                
                r_data[38115] <= r_data[38114];
                
                r_data[38116] <= r_data[38115];
                
                r_data[38117] <= r_data[38116];
                
                r_data[38118] <= r_data[38117];
                
                r_data[38119] <= r_data[38118];
                
                r_data[38120] <= r_data[38119];
                
                r_data[38121] <= r_data[38120];
                
                r_data[38122] <= r_data[38121];
                
                r_data[38123] <= r_data[38122];
                
                r_data[38124] <= r_data[38123];
                
                r_data[38125] <= r_data[38124];
                
                r_data[38126] <= r_data[38125];
                
                r_data[38127] <= r_data[38126];
                
                r_data[38128] <= r_data[38127];
                
                r_data[38129] <= r_data[38128];
                
                r_data[38130] <= r_data[38129];
                
                r_data[38131] <= r_data[38130];
                
                r_data[38132] <= r_data[38131];
                
                r_data[38133] <= r_data[38132];
                
                r_data[38134] <= r_data[38133];
                
                r_data[38135] <= r_data[38134];
                
                r_data[38136] <= r_data[38135];
                
                r_data[38137] <= r_data[38136];
                
                r_data[38138] <= r_data[38137];
                
                r_data[38139] <= r_data[38138];
                
                r_data[38140] <= r_data[38139];
                
                r_data[38141] <= r_data[38140];
                
                r_data[38142] <= r_data[38141];
                
                r_data[38143] <= r_data[38142];
                
                r_data[38144] <= r_data[38143];
                
                r_data[38145] <= r_data[38144];
                
                r_data[38146] <= r_data[38145];
                
                r_data[38147] <= r_data[38146];
                
                r_data[38148] <= r_data[38147];
                
                r_data[38149] <= r_data[38148];
                
                r_data[38150] <= r_data[38149];
                
                r_data[38151] <= r_data[38150];
                
                r_data[38152] <= r_data[38151];
                
                r_data[38153] <= r_data[38152];
                
                r_data[38154] <= r_data[38153];
                
                r_data[38155] <= r_data[38154];
                
                r_data[38156] <= r_data[38155];
                
                r_data[38157] <= r_data[38156];
                
                r_data[38158] <= r_data[38157];
                
                r_data[38159] <= r_data[38158];
                
                r_data[38160] <= r_data[38159];
                
                r_data[38161] <= r_data[38160];
                
                r_data[38162] <= r_data[38161];
                
                r_data[38163] <= r_data[38162];
                
                r_data[38164] <= r_data[38163];
                
                r_data[38165] <= r_data[38164];
                
                r_data[38166] <= r_data[38165];
                
                r_data[38167] <= r_data[38166];
                
                r_data[38168] <= r_data[38167];
                
                r_data[38169] <= r_data[38168];
                
                r_data[38170] <= r_data[38169];
                
                r_data[38171] <= r_data[38170];
                
                r_data[38172] <= r_data[38171];
                
                r_data[38173] <= r_data[38172];
                
                r_data[38174] <= r_data[38173];
                
                r_data[38175] <= r_data[38174];
                
                r_data[38176] <= r_data[38175];
                
                r_data[38177] <= r_data[38176];
                
                r_data[38178] <= r_data[38177];
                
                r_data[38179] <= r_data[38178];
                
                r_data[38180] <= r_data[38179];
                
                r_data[38181] <= r_data[38180];
                
                r_data[38182] <= r_data[38181];
                
                r_data[38183] <= r_data[38182];
                
                r_data[38184] <= r_data[38183];
                
                r_data[38185] <= r_data[38184];
                
                r_data[38186] <= r_data[38185];
                
                r_data[38187] <= r_data[38186];
                
                r_data[38188] <= r_data[38187];
                
                r_data[38189] <= r_data[38188];
                
                r_data[38190] <= r_data[38189];
                
                r_data[38191] <= r_data[38190];
                
                r_data[38192] <= r_data[38191];
                
                r_data[38193] <= r_data[38192];
                
                r_data[38194] <= r_data[38193];
                
                r_data[38195] <= r_data[38194];
                
                r_data[38196] <= r_data[38195];
                
                r_data[38197] <= r_data[38196];
                
                r_data[38198] <= r_data[38197];
                
                r_data[38199] <= r_data[38198];
                
                r_data[38200] <= r_data[38199];
                
                r_data[38201] <= r_data[38200];
                
                r_data[38202] <= r_data[38201];
                
                r_data[38203] <= r_data[38202];
                
                r_data[38204] <= r_data[38203];
                
                r_data[38205] <= r_data[38204];
                
                r_data[38206] <= r_data[38205];
                
                r_data[38207] <= r_data[38206];
                
                r_data[38208] <= r_data[38207];
                
                r_data[38209] <= r_data[38208];
                
                r_data[38210] <= r_data[38209];
                
                r_data[38211] <= r_data[38210];
                
                r_data[38212] <= r_data[38211];
                
                r_data[38213] <= r_data[38212];
                
                r_data[38214] <= r_data[38213];
                
                r_data[38215] <= r_data[38214];
                
                r_data[38216] <= r_data[38215];
                
                r_data[38217] <= r_data[38216];
                
                r_data[38218] <= r_data[38217];
                
                r_data[38219] <= r_data[38218];
                
                r_data[38220] <= r_data[38219];
                
                r_data[38221] <= r_data[38220];
                
                r_data[38222] <= r_data[38221];
                
                r_data[38223] <= r_data[38222];
                
                r_data[38224] <= r_data[38223];
                
                r_data[38225] <= r_data[38224];
                
                r_data[38226] <= r_data[38225];
                
                r_data[38227] <= r_data[38226];
                
                r_data[38228] <= r_data[38227];
                
                r_data[38229] <= r_data[38228];
                
                r_data[38230] <= r_data[38229];
                
                r_data[38231] <= r_data[38230];
                
                r_data[38232] <= r_data[38231];
                
                r_data[38233] <= r_data[38232];
                
                r_data[38234] <= r_data[38233];
                
                r_data[38235] <= r_data[38234];
                
                r_data[38236] <= r_data[38235];
                
                r_data[38237] <= r_data[38236];
                
                r_data[38238] <= r_data[38237];
                
                r_data[38239] <= r_data[38238];
                
                r_data[38240] <= r_data[38239];
                
                r_data[38241] <= r_data[38240];
                
                r_data[38242] <= r_data[38241];
                
                r_data[38243] <= r_data[38242];
                
                r_data[38244] <= r_data[38243];
                
                r_data[38245] <= r_data[38244];
                
                r_data[38246] <= r_data[38245];
                
                r_data[38247] <= r_data[38246];
                
                r_data[38248] <= r_data[38247];
                
                r_data[38249] <= r_data[38248];
                
                r_data[38250] <= r_data[38249];
                
                r_data[38251] <= r_data[38250];
                
                r_data[38252] <= r_data[38251];
                
                r_data[38253] <= r_data[38252];
                
                r_data[38254] <= r_data[38253];
                
                r_data[38255] <= r_data[38254];
                
                r_data[38256] <= r_data[38255];
                
                r_data[38257] <= r_data[38256];
                
                r_data[38258] <= r_data[38257];
                
                r_data[38259] <= r_data[38258];
                
                r_data[38260] <= r_data[38259];
                
                r_data[38261] <= r_data[38260];
                
                r_data[38262] <= r_data[38261];
                
                r_data[38263] <= r_data[38262];
                
                r_data[38264] <= r_data[38263];
                
                r_data[38265] <= r_data[38264];
                
                r_data[38266] <= r_data[38265];
                
                r_data[38267] <= r_data[38266];
                
                r_data[38268] <= r_data[38267];
                
                r_data[38269] <= r_data[38268];
                
                r_data[38270] <= r_data[38269];
                
                r_data[38271] <= r_data[38270];
                
                r_data[38272] <= r_data[38271];
                
                r_data[38273] <= r_data[38272];
                
                r_data[38274] <= r_data[38273];
                
                r_data[38275] <= r_data[38274];
                
                r_data[38276] <= r_data[38275];
                
                r_data[38277] <= r_data[38276];
                
                r_data[38278] <= r_data[38277];
                
                r_data[38279] <= r_data[38278];
                
                r_data[38280] <= r_data[38279];
                
                r_data[38281] <= r_data[38280];
                
                r_data[38282] <= r_data[38281];
                
                r_data[38283] <= r_data[38282];
                
                r_data[38284] <= r_data[38283];
                
                r_data[38285] <= r_data[38284];
                
                r_data[38286] <= r_data[38285];
                
                r_data[38287] <= r_data[38286];
                
                r_data[38288] <= r_data[38287];
                
                r_data[38289] <= r_data[38288];
                
                r_data[38290] <= r_data[38289];
                
                r_data[38291] <= r_data[38290];
                
                r_data[38292] <= r_data[38291];
                
                r_data[38293] <= r_data[38292];
                
                r_data[38294] <= r_data[38293];
                
                r_data[38295] <= r_data[38294];
                
                r_data[38296] <= r_data[38295];
                
                r_data[38297] <= r_data[38296];
                
                r_data[38298] <= r_data[38297];
                
                r_data[38299] <= r_data[38298];
                
                r_data[38300] <= r_data[38299];
                
                r_data[38301] <= r_data[38300];
                
                r_data[38302] <= r_data[38301];
                
                r_data[38303] <= r_data[38302];
                
                r_data[38304] <= r_data[38303];
                
                r_data[38305] <= r_data[38304];
                
                r_data[38306] <= r_data[38305];
                
                r_data[38307] <= r_data[38306];
                
                r_data[38308] <= r_data[38307];
                
                r_data[38309] <= r_data[38308];
                
                r_data[38310] <= r_data[38309];
                
                r_data[38311] <= r_data[38310];
                
                r_data[38312] <= r_data[38311];
                
                r_data[38313] <= r_data[38312];
                
                r_data[38314] <= r_data[38313];
                
                r_data[38315] <= r_data[38314];
                
                r_data[38316] <= r_data[38315];
                
                r_data[38317] <= r_data[38316];
                
                r_data[38318] <= r_data[38317];
                
                r_data[38319] <= r_data[38318];
                
                r_data[38320] <= r_data[38319];
                
                r_data[38321] <= r_data[38320];
                
                r_data[38322] <= r_data[38321];
                
                r_data[38323] <= r_data[38322];
                
                r_data[38324] <= r_data[38323];
                
                r_data[38325] <= r_data[38324];
                
                r_data[38326] <= r_data[38325];
                
                r_data[38327] <= r_data[38326];
                
                r_data[38328] <= r_data[38327];
                
                r_data[38329] <= r_data[38328];
                
                r_data[38330] <= r_data[38329];
                
                r_data[38331] <= r_data[38330];
                
                r_data[38332] <= r_data[38331];
                
                r_data[38333] <= r_data[38332];
                
                r_data[38334] <= r_data[38333];
                
                r_data[38335] <= r_data[38334];
                
                r_data[38336] <= r_data[38335];
                
                r_data[38337] <= r_data[38336];
                
                r_data[38338] <= r_data[38337];
                
                r_data[38339] <= r_data[38338];
                
                r_data[38340] <= r_data[38339];
                
                r_data[38341] <= r_data[38340];
                
                r_data[38342] <= r_data[38341];
                
                r_data[38343] <= r_data[38342];
                
                r_data[38344] <= r_data[38343];
                
                r_data[38345] <= r_data[38344];
                
                r_data[38346] <= r_data[38345];
                
                r_data[38347] <= r_data[38346];
                
                r_data[38348] <= r_data[38347];
                
                r_data[38349] <= r_data[38348];
                
                r_data[38350] <= r_data[38349];
                
                r_data[38351] <= r_data[38350];
                
                r_data[38352] <= r_data[38351];
                
                r_data[38353] <= r_data[38352];
                
                r_data[38354] <= r_data[38353];
                
                r_data[38355] <= r_data[38354];
                
                r_data[38356] <= r_data[38355];
                
                r_data[38357] <= r_data[38356];
                
                r_data[38358] <= r_data[38357];
                
                r_data[38359] <= r_data[38358];
                
                r_data[38360] <= r_data[38359];
                
                r_data[38361] <= r_data[38360];
                
                r_data[38362] <= r_data[38361];
                
                r_data[38363] <= r_data[38362];
                
                r_data[38364] <= r_data[38363];
                
                r_data[38365] <= r_data[38364];
                
                r_data[38366] <= r_data[38365];
                
                r_data[38367] <= r_data[38366];
                
                r_data[38368] <= r_data[38367];
                
                r_data[38369] <= r_data[38368];
                
                r_data[38370] <= r_data[38369];
                
                r_data[38371] <= r_data[38370];
                
                r_data[38372] <= r_data[38371];
                
                r_data[38373] <= r_data[38372];
                
                r_data[38374] <= r_data[38373];
                
                r_data[38375] <= r_data[38374];
                
                r_data[38376] <= r_data[38375];
                
                r_data[38377] <= r_data[38376];
                
                r_data[38378] <= r_data[38377];
                
                r_data[38379] <= r_data[38378];
                
                r_data[38380] <= r_data[38379];
                
                r_data[38381] <= r_data[38380];
                
                r_data[38382] <= r_data[38381];
                
                r_data[38383] <= r_data[38382];
                
                r_data[38384] <= r_data[38383];
                
                r_data[38385] <= r_data[38384];
                
                r_data[38386] <= r_data[38385];
                
                r_data[38387] <= r_data[38386];
                
                r_data[38388] <= r_data[38387];
                
                r_data[38389] <= r_data[38388];
                
                r_data[38390] <= r_data[38389];
                
                r_data[38391] <= r_data[38390];
                
                r_data[38392] <= r_data[38391];
                
                r_data[38393] <= r_data[38392];
                
                r_data[38394] <= r_data[38393];
                
                r_data[38395] <= r_data[38394];
                
                r_data[38396] <= r_data[38395];
                
                r_data[38397] <= r_data[38396];
                
                r_data[38398] <= r_data[38397];
                
                r_data[38399] <= r_data[38398];
                
                r_data[38400] <= r_data[38399];
                
                r_data[38401] <= r_data[38400];
                
                r_data[38402] <= r_data[38401];
                
                r_data[38403] <= r_data[38402];
                
                r_data[38404] <= r_data[38403];
                
                r_data[38405] <= r_data[38404];
                
                r_data[38406] <= r_data[38405];
                
                r_data[38407] <= r_data[38406];
                
                r_data[38408] <= r_data[38407];
                
                r_data[38409] <= r_data[38408];
                
                r_data[38410] <= r_data[38409];
                
                r_data[38411] <= r_data[38410];
                
                r_data[38412] <= r_data[38411];
                
                r_data[38413] <= r_data[38412];
                
                r_data[38414] <= r_data[38413];
                
                r_data[38415] <= r_data[38414];
                
                r_data[38416] <= r_data[38415];
                
                r_data[38417] <= r_data[38416];
                
                r_data[38418] <= r_data[38417];
                
                r_data[38419] <= r_data[38418];
                
                r_data[38420] <= r_data[38419];
                
                r_data[38421] <= r_data[38420];
                
                r_data[38422] <= r_data[38421];
                
                r_data[38423] <= r_data[38422];
                
                r_data[38424] <= r_data[38423];
                
                r_data[38425] <= r_data[38424];
                
                r_data[38426] <= r_data[38425];
                
                r_data[38427] <= r_data[38426];
                
                r_data[38428] <= r_data[38427];
                
                r_data[38429] <= r_data[38428];
                
                r_data[38430] <= r_data[38429];
                
                r_data[38431] <= r_data[38430];
                
                r_data[38432] <= r_data[38431];
                
                r_data[38433] <= r_data[38432];
                
                r_data[38434] <= r_data[38433];
                
                r_data[38435] <= r_data[38434];
                
                r_data[38436] <= r_data[38435];
                
                r_data[38437] <= r_data[38436];
                
                r_data[38438] <= r_data[38437];
                
                r_data[38439] <= r_data[38438];
                
                r_data[38440] <= r_data[38439];
                
                r_data[38441] <= r_data[38440];
                
                r_data[38442] <= r_data[38441];
                
                r_data[38443] <= r_data[38442];
                
                r_data[38444] <= r_data[38443];
                
                r_data[38445] <= r_data[38444];
                
                r_data[38446] <= r_data[38445];
                
                r_data[38447] <= r_data[38446];
                
                r_data[38448] <= r_data[38447];
                
                r_data[38449] <= r_data[38448];
                
                r_data[38450] <= r_data[38449];
                
                r_data[38451] <= r_data[38450];
                
                r_data[38452] <= r_data[38451];
                
                r_data[38453] <= r_data[38452];
                
                r_data[38454] <= r_data[38453];
                
                r_data[38455] <= r_data[38454];
                
                r_data[38456] <= r_data[38455];
                
                r_data[38457] <= r_data[38456];
                
                r_data[38458] <= r_data[38457];
                
                r_data[38459] <= r_data[38458];
                
                r_data[38460] <= r_data[38459];
                
                r_data[38461] <= r_data[38460];
                
                r_data[38462] <= r_data[38461];
                
                r_data[38463] <= r_data[38462];
                
                r_data[38464] <= r_data[38463];
                
                r_data[38465] <= r_data[38464];
                
                r_data[38466] <= r_data[38465];
                
                r_data[38467] <= r_data[38466];
                
                r_data[38468] <= r_data[38467];
                
                r_data[38469] <= r_data[38468];
                
                r_data[38470] <= r_data[38469];
                
                r_data[38471] <= r_data[38470];
                
                r_data[38472] <= r_data[38471];
                
                r_data[38473] <= r_data[38472];
                
                r_data[38474] <= r_data[38473];
                
                r_data[38475] <= r_data[38474];
                
                r_data[38476] <= r_data[38475];
                
                r_data[38477] <= r_data[38476];
                
                r_data[38478] <= r_data[38477];
                
                r_data[38479] <= r_data[38478];
                
                r_data[38480] <= r_data[38479];
                
                r_data[38481] <= r_data[38480];
                
                r_data[38482] <= r_data[38481];
                
                r_data[38483] <= r_data[38482];
                
                r_data[38484] <= r_data[38483];
                
                r_data[38485] <= r_data[38484];
                
                r_data[38486] <= r_data[38485];
                
                r_data[38487] <= r_data[38486];
                
                r_data[38488] <= r_data[38487];
                
                r_data[38489] <= r_data[38488];
                
                r_data[38490] <= r_data[38489];
                
                r_data[38491] <= r_data[38490];
                
                r_data[38492] <= r_data[38491];
                
                r_data[38493] <= r_data[38492];
                
                r_data[38494] <= r_data[38493];
                
                r_data[38495] <= r_data[38494];
                
                r_data[38496] <= r_data[38495];
                
                r_data[38497] <= r_data[38496];
                
                r_data[38498] <= r_data[38497];
                
                r_data[38499] <= r_data[38498];
                
                r_data[38500] <= r_data[38499];
                
                r_data[38501] <= r_data[38500];
                
                r_data[38502] <= r_data[38501];
                
                r_data[38503] <= r_data[38502];
                
                r_data[38504] <= r_data[38503];
                
                r_data[38505] <= r_data[38504];
                
                r_data[38506] <= r_data[38505];
                
                r_data[38507] <= r_data[38506];
                
                r_data[38508] <= r_data[38507];
                
                r_data[38509] <= r_data[38508];
                
                r_data[38510] <= r_data[38509];
                
                r_data[38511] <= r_data[38510];
                
                r_data[38512] <= r_data[38511];
                
                r_data[38513] <= r_data[38512];
                
                r_data[38514] <= r_data[38513];
                
                r_data[38515] <= r_data[38514];
                
                r_data[38516] <= r_data[38515];
                
                r_data[38517] <= r_data[38516];
                
                r_data[38518] <= r_data[38517];
                
                r_data[38519] <= r_data[38518];
                
                r_data[38520] <= r_data[38519];
                
                r_data[38521] <= r_data[38520];
                
                r_data[38522] <= r_data[38521];
                
                r_data[38523] <= r_data[38522];
                
                r_data[38524] <= r_data[38523];
                
                r_data[38525] <= r_data[38524];
                
                r_data[38526] <= r_data[38525];
                
                r_data[38527] <= r_data[38526];
                
                r_data[38528] <= r_data[38527];
                
                r_data[38529] <= r_data[38528];
                
                r_data[38530] <= r_data[38529];
                
                r_data[38531] <= r_data[38530];
                
                r_data[38532] <= r_data[38531];
                
                r_data[38533] <= r_data[38532];
                
                r_data[38534] <= r_data[38533];
                
                r_data[38535] <= r_data[38534];
                
                r_data[38536] <= r_data[38535];
                
                r_data[38537] <= r_data[38536];
                
                r_data[38538] <= r_data[38537];
                
                r_data[38539] <= r_data[38538];
                
                r_data[38540] <= r_data[38539];
                
                r_data[38541] <= r_data[38540];
                
                r_data[38542] <= r_data[38541];
                
                r_data[38543] <= r_data[38542];
                
                r_data[38544] <= r_data[38543];
                
                r_data[38545] <= r_data[38544];
                
                r_data[38546] <= r_data[38545];
                
                r_data[38547] <= r_data[38546];
                
                r_data[38548] <= r_data[38547];
                
                r_data[38549] <= r_data[38548];
                
                r_data[38550] <= r_data[38549];
                
                r_data[38551] <= r_data[38550];
                
                r_data[38552] <= r_data[38551];
                
                r_data[38553] <= r_data[38552];
                
                r_data[38554] <= r_data[38553];
                
                r_data[38555] <= r_data[38554];
                
                r_data[38556] <= r_data[38555];
                
                r_data[38557] <= r_data[38556];
                
                r_data[38558] <= r_data[38557];
                
                r_data[38559] <= r_data[38558];
                
                r_data[38560] <= r_data[38559];
                
                r_data[38561] <= r_data[38560];
                
                r_data[38562] <= r_data[38561];
                
                r_data[38563] <= r_data[38562];
                
                r_data[38564] <= r_data[38563];
                
                r_data[38565] <= r_data[38564];
                
                r_data[38566] <= r_data[38565];
                
                r_data[38567] <= r_data[38566];
                
                r_data[38568] <= r_data[38567];
                
                r_data[38569] <= r_data[38568];
                
                r_data[38570] <= r_data[38569];
                
                r_data[38571] <= r_data[38570];
                
                r_data[38572] <= r_data[38571];
                
                r_data[38573] <= r_data[38572];
                
                r_data[38574] <= r_data[38573];
                
                r_data[38575] <= r_data[38574];
                
                r_data[38576] <= r_data[38575];
                
                r_data[38577] <= r_data[38576];
                
                r_data[38578] <= r_data[38577];
                
                r_data[38579] <= r_data[38578];
                
                r_data[38580] <= r_data[38579];
                
                r_data[38581] <= r_data[38580];
                
                r_data[38582] <= r_data[38581];
                
                r_data[38583] <= r_data[38582];
                
                r_data[38584] <= r_data[38583];
                
                r_data[38585] <= r_data[38584];
                
                r_data[38586] <= r_data[38585];
                
                r_data[38587] <= r_data[38586];
                
                r_data[38588] <= r_data[38587];
                
                r_data[38589] <= r_data[38588];
                
                r_data[38590] <= r_data[38589];
                
                r_data[38591] <= r_data[38590];
                
                r_data[38592] <= r_data[38591];
                
                r_data[38593] <= r_data[38592];
                
                r_data[38594] <= r_data[38593];
                
                r_data[38595] <= r_data[38594];
                
                r_data[38596] <= r_data[38595];
                
                r_data[38597] <= r_data[38596];
                
                r_data[38598] <= r_data[38597];
                
                r_data[38599] <= r_data[38598];
                
                r_data[38600] <= r_data[38599];
                
                r_data[38601] <= r_data[38600];
                
                r_data[38602] <= r_data[38601];
                
                r_data[38603] <= r_data[38602];
                
                r_data[38604] <= r_data[38603];
                
                r_data[38605] <= r_data[38604];
                
                r_data[38606] <= r_data[38605];
                
                r_data[38607] <= r_data[38606];
                
                r_data[38608] <= r_data[38607];
                
                r_data[38609] <= r_data[38608];
                
                r_data[38610] <= r_data[38609];
                
                r_data[38611] <= r_data[38610];
                
                r_data[38612] <= r_data[38611];
                
                r_data[38613] <= r_data[38612];
                
                r_data[38614] <= r_data[38613];
                
                r_data[38615] <= r_data[38614];
                
                r_data[38616] <= r_data[38615];
                
                r_data[38617] <= r_data[38616];
                
                r_data[38618] <= r_data[38617];
                
                r_data[38619] <= r_data[38618];
                
                r_data[38620] <= r_data[38619];
                
                r_data[38621] <= r_data[38620];
                
                r_data[38622] <= r_data[38621];
                
                r_data[38623] <= r_data[38622];
                
                r_data[38624] <= r_data[38623];
                
                r_data[38625] <= r_data[38624];
                
                r_data[38626] <= r_data[38625];
                
                r_data[38627] <= r_data[38626];
                
                r_data[38628] <= r_data[38627];
                
                r_data[38629] <= r_data[38628];
                
                r_data[38630] <= r_data[38629];
                
                r_data[38631] <= r_data[38630];
                
                r_data[38632] <= r_data[38631];
                
                r_data[38633] <= r_data[38632];
                
                r_data[38634] <= r_data[38633];
                
                r_data[38635] <= r_data[38634];
                
                r_data[38636] <= r_data[38635];
                
                r_data[38637] <= r_data[38636];
                
                r_data[38638] <= r_data[38637];
                
                r_data[38639] <= r_data[38638];
                
                r_data[38640] <= r_data[38639];
                
                r_data[38641] <= r_data[38640];
                
                r_data[38642] <= r_data[38641];
                
                r_data[38643] <= r_data[38642];
                
                r_data[38644] <= r_data[38643];
                
                r_data[38645] <= r_data[38644];
                
                r_data[38646] <= r_data[38645];
                
                r_data[38647] <= r_data[38646];
                
                r_data[38648] <= r_data[38647];
                
                r_data[38649] <= r_data[38648];
                
                r_data[38650] <= r_data[38649];
                
                r_data[38651] <= r_data[38650];
                
                r_data[38652] <= r_data[38651];
                
                r_data[38653] <= r_data[38652];
                
                r_data[38654] <= r_data[38653];
                
                r_data[38655] <= r_data[38654];
                
                r_data[38656] <= r_data[38655];
                
                r_data[38657] <= r_data[38656];
                
                r_data[38658] <= r_data[38657];
                
                r_data[38659] <= r_data[38658];
                
                r_data[38660] <= r_data[38659];
                
                r_data[38661] <= r_data[38660];
                
                r_data[38662] <= r_data[38661];
                
                r_data[38663] <= r_data[38662];
                
                r_data[38664] <= r_data[38663];
                
                r_data[38665] <= r_data[38664];
                
                r_data[38666] <= r_data[38665];
                
                r_data[38667] <= r_data[38666];
                
                r_data[38668] <= r_data[38667];
                
                r_data[38669] <= r_data[38668];
                
                r_data[38670] <= r_data[38669];
                
                r_data[38671] <= r_data[38670];
                
                r_data[38672] <= r_data[38671];
                
                r_data[38673] <= r_data[38672];
                
                r_data[38674] <= r_data[38673];
                
                r_data[38675] <= r_data[38674];
                
                r_data[38676] <= r_data[38675];
                
                r_data[38677] <= r_data[38676];
                
                r_data[38678] <= r_data[38677];
                
                r_data[38679] <= r_data[38678];
                
                r_data[38680] <= r_data[38679];
                
                r_data[38681] <= r_data[38680];
                
                r_data[38682] <= r_data[38681];
                
                r_data[38683] <= r_data[38682];
                
                r_data[38684] <= r_data[38683];
                
                r_data[38685] <= r_data[38684];
                
                r_data[38686] <= r_data[38685];
                
                r_data[38687] <= r_data[38686];
                
                r_data[38688] <= r_data[38687];
                
                r_data[38689] <= r_data[38688];
                
                r_data[38690] <= r_data[38689];
                
                r_data[38691] <= r_data[38690];
                
                r_data[38692] <= r_data[38691];
                
                r_data[38693] <= r_data[38692];
                
                r_data[38694] <= r_data[38693];
                
                r_data[38695] <= r_data[38694];
                
                r_data[38696] <= r_data[38695];
                
                r_data[38697] <= r_data[38696];
                
                r_data[38698] <= r_data[38697];
                
                r_data[38699] <= r_data[38698];
                
                r_data[38700] <= r_data[38699];
                
                r_data[38701] <= r_data[38700];
                
                r_data[38702] <= r_data[38701];
                
                r_data[38703] <= r_data[38702];
                
                r_data[38704] <= r_data[38703];
                
                r_data[38705] <= r_data[38704];
                
                r_data[38706] <= r_data[38705];
                
                r_data[38707] <= r_data[38706];
                
                r_data[38708] <= r_data[38707];
                
                r_data[38709] <= r_data[38708];
                
                r_data[38710] <= r_data[38709];
                
                r_data[38711] <= r_data[38710];
                
                r_data[38712] <= r_data[38711];
                
                r_data[38713] <= r_data[38712];
                
                r_data[38714] <= r_data[38713];
                
                r_data[38715] <= r_data[38714];
                
                r_data[38716] <= r_data[38715];
                
                r_data[38717] <= r_data[38716];
                
                r_data[38718] <= r_data[38717];
                
                r_data[38719] <= r_data[38718];
                
                r_data[38720] <= r_data[38719];
                
                r_data[38721] <= r_data[38720];
                
                r_data[38722] <= r_data[38721];
                
                r_data[38723] <= r_data[38722];
                
                r_data[38724] <= r_data[38723];
                
                r_data[38725] <= r_data[38724];
                
                r_data[38726] <= r_data[38725];
                
                r_data[38727] <= r_data[38726];
                
                r_data[38728] <= r_data[38727];
                
                r_data[38729] <= r_data[38728];
                
                r_data[38730] <= r_data[38729];
                
                r_data[38731] <= r_data[38730];
                
                r_data[38732] <= r_data[38731];
                
                r_data[38733] <= r_data[38732];
                
                r_data[38734] <= r_data[38733];
                
                r_data[38735] <= r_data[38734];
                
                r_data[38736] <= r_data[38735];
                
                r_data[38737] <= r_data[38736];
                
                r_data[38738] <= r_data[38737];
                
                r_data[38739] <= r_data[38738];
                
                r_data[38740] <= r_data[38739];
                
                r_data[38741] <= r_data[38740];
                
                r_data[38742] <= r_data[38741];
                
                r_data[38743] <= r_data[38742];
                
                r_data[38744] <= r_data[38743];
                
                r_data[38745] <= r_data[38744];
                
                r_data[38746] <= r_data[38745];
                
                r_data[38747] <= r_data[38746];
                
                r_data[38748] <= r_data[38747];
                
                r_data[38749] <= r_data[38748];
                
                r_data[38750] <= r_data[38749];
                
                r_data[38751] <= r_data[38750];
                
                r_data[38752] <= r_data[38751];
                
                r_data[38753] <= r_data[38752];
                
                r_data[38754] <= r_data[38753];
                
                r_data[38755] <= r_data[38754];
                
                r_data[38756] <= r_data[38755];
                
                r_data[38757] <= r_data[38756];
                
                r_data[38758] <= r_data[38757];
                
                r_data[38759] <= r_data[38758];
                
                r_data[38760] <= r_data[38759];
                
                r_data[38761] <= r_data[38760];
                
                r_data[38762] <= r_data[38761];
                
                r_data[38763] <= r_data[38762];
                
                r_data[38764] <= r_data[38763];
                
                r_data[38765] <= r_data[38764];
                
                r_data[38766] <= r_data[38765];
                
                r_data[38767] <= r_data[38766];
                
                r_data[38768] <= r_data[38767];
                
                r_data[38769] <= r_data[38768];
                
                r_data[38770] <= r_data[38769];
                
                r_data[38771] <= r_data[38770];
                
                r_data[38772] <= r_data[38771];
                
                r_data[38773] <= r_data[38772];
                
                r_data[38774] <= r_data[38773];
                
                r_data[38775] <= r_data[38774];
                
                r_data[38776] <= r_data[38775];
                
                r_data[38777] <= r_data[38776];
                
                r_data[38778] <= r_data[38777];
                
                r_data[38779] <= r_data[38778];
                
                r_data[38780] <= r_data[38779];
                
                r_data[38781] <= r_data[38780];
                
                r_data[38782] <= r_data[38781];
                
                r_data[38783] <= r_data[38782];
                
                r_data[38784] <= r_data[38783];
                
                r_data[38785] <= r_data[38784];
                
                r_data[38786] <= r_data[38785];
                
                r_data[38787] <= r_data[38786];
                
                r_data[38788] <= r_data[38787];
                
                r_data[38789] <= r_data[38788];
                
                r_data[38790] <= r_data[38789];
                
                r_data[38791] <= r_data[38790];
                
                r_data[38792] <= r_data[38791];
                
                r_data[38793] <= r_data[38792];
                
                r_data[38794] <= r_data[38793];
                
                r_data[38795] <= r_data[38794];
                
                r_data[38796] <= r_data[38795];
                
                r_data[38797] <= r_data[38796];
                
                r_data[38798] <= r_data[38797];
                
                r_data[38799] <= r_data[38798];
                
                r_data[38800] <= r_data[38799];
                
                r_data[38801] <= r_data[38800];
                
                r_data[38802] <= r_data[38801];
                
                r_data[38803] <= r_data[38802];
                
                r_data[38804] <= r_data[38803];
                
                r_data[38805] <= r_data[38804];
                
                r_data[38806] <= r_data[38805];
                
                r_data[38807] <= r_data[38806];
                
                r_data[38808] <= r_data[38807];
                
                r_data[38809] <= r_data[38808];
                
                r_data[38810] <= r_data[38809];
                
                r_data[38811] <= r_data[38810];
                
                r_data[38812] <= r_data[38811];
                
                r_data[38813] <= r_data[38812];
                
                r_data[38814] <= r_data[38813];
                
                r_data[38815] <= r_data[38814];
                
                r_data[38816] <= r_data[38815];
                
                r_data[38817] <= r_data[38816];
                
                r_data[38818] <= r_data[38817];
                
                r_data[38819] <= r_data[38818];
                
                r_data[38820] <= r_data[38819];
                
                r_data[38821] <= r_data[38820];
                
                r_data[38822] <= r_data[38821];
                
                r_data[38823] <= r_data[38822];
                
                r_data[38824] <= r_data[38823];
                
                r_data[38825] <= r_data[38824];
                
                r_data[38826] <= r_data[38825];
                
                r_data[38827] <= r_data[38826];
                
                r_data[38828] <= r_data[38827];
                
                r_data[38829] <= r_data[38828];
                
                r_data[38830] <= r_data[38829];
                
                r_data[38831] <= r_data[38830];
                
                r_data[38832] <= r_data[38831];
                
                r_data[38833] <= r_data[38832];
                
                r_data[38834] <= r_data[38833];
                
                r_data[38835] <= r_data[38834];
                
                r_data[38836] <= r_data[38835];
                
                r_data[38837] <= r_data[38836];
                
                r_data[38838] <= r_data[38837];
                
                r_data[38839] <= r_data[38838];
                
                r_data[38840] <= r_data[38839];
                
                r_data[38841] <= r_data[38840];
                
                r_data[38842] <= r_data[38841];
                
                r_data[38843] <= r_data[38842];
                
                r_data[38844] <= r_data[38843];
                
                r_data[38845] <= r_data[38844];
                
                r_data[38846] <= r_data[38845];
                
                r_data[38847] <= r_data[38846];
                
                r_data[38848] <= r_data[38847];
                
                r_data[38849] <= r_data[38848];
                
                r_data[38850] <= r_data[38849];
                
                r_data[38851] <= r_data[38850];
                
                r_data[38852] <= r_data[38851];
                
                r_data[38853] <= r_data[38852];
                
                r_data[38854] <= r_data[38853];
                
                r_data[38855] <= r_data[38854];
                
                r_data[38856] <= r_data[38855];
                
                r_data[38857] <= r_data[38856];
                
                r_data[38858] <= r_data[38857];
                
                r_data[38859] <= r_data[38858];
                
                r_data[38860] <= r_data[38859];
                
                r_data[38861] <= r_data[38860];
                
                r_data[38862] <= r_data[38861];
                
                r_data[38863] <= r_data[38862];
                
                r_data[38864] <= r_data[38863];
                
                r_data[38865] <= r_data[38864];
                
                r_data[38866] <= r_data[38865];
                
                r_data[38867] <= r_data[38866];
                
                r_data[38868] <= r_data[38867];
                
                r_data[38869] <= r_data[38868];
                
                r_data[38870] <= r_data[38869];
                
                r_data[38871] <= r_data[38870];
                
                r_data[38872] <= r_data[38871];
                
                r_data[38873] <= r_data[38872];
                
                r_data[38874] <= r_data[38873];
                
                r_data[38875] <= r_data[38874];
                
                r_data[38876] <= r_data[38875];
                
                r_data[38877] <= r_data[38876];
                
                r_data[38878] <= r_data[38877];
                
                r_data[38879] <= r_data[38878];
                
                r_data[38880] <= r_data[38879];
                
                r_data[38881] <= r_data[38880];
                
                r_data[38882] <= r_data[38881];
                
                r_data[38883] <= r_data[38882];
                
                r_data[38884] <= r_data[38883];
                
                r_data[38885] <= r_data[38884];
                
                r_data[38886] <= r_data[38885];
                
                r_data[38887] <= r_data[38886];
                
                r_data[38888] <= r_data[38887];
                
                r_data[38889] <= r_data[38888];
                
                r_data[38890] <= r_data[38889];
                
                r_data[38891] <= r_data[38890];
                
                r_data[38892] <= r_data[38891];
                
                r_data[38893] <= r_data[38892];
                
                r_data[38894] <= r_data[38893];
                
                r_data[38895] <= r_data[38894];
                
                r_data[38896] <= r_data[38895];
                
                r_data[38897] <= r_data[38896];
                
                r_data[38898] <= r_data[38897];
                
                r_data[38899] <= r_data[38898];
                
                r_data[38900] <= r_data[38899];
                
                r_data[38901] <= r_data[38900];
                
                r_data[38902] <= r_data[38901];
                
                r_data[38903] <= r_data[38902];
                
                r_data[38904] <= r_data[38903];
                
                r_data[38905] <= r_data[38904];
                
                r_data[38906] <= r_data[38905];
                
                r_data[38907] <= r_data[38906];
                
                r_data[38908] <= r_data[38907];
                
                r_data[38909] <= r_data[38908];
                
                r_data[38910] <= r_data[38909];
                
                r_data[38911] <= r_data[38910];
                
                r_data[38912] <= r_data[38911];
                
                r_data[38913] <= r_data[38912];
                
                r_data[38914] <= r_data[38913];
                
                r_data[38915] <= r_data[38914];
                
                r_data[38916] <= r_data[38915];
                
                r_data[38917] <= r_data[38916];
                
                r_data[38918] <= r_data[38917];
                
                r_data[38919] <= r_data[38918];
                
                r_data[38920] <= r_data[38919];
                
                r_data[38921] <= r_data[38920];
                
                r_data[38922] <= r_data[38921];
                
                r_data[38923] <= r_data[38922];
                
                r_data[38924] <= r_data[38923];
                
                r_data[38925] <= r_data[38924];
                
                r_data[38926] <= r_data[38925];
                
                r_data[38927] <= r_data[38926];
                
                r_data[38928] <= r_data[38927];
                
                r_data[38929] <= r_data[38928];
                
                r_data[38930] <= r_data[38929];
                
                r_data[38931] <= r_data[38930];
                
                r_data[38932] <= r_data[38931];
                
                r_data[38933] <= r_data[38932];
                
                r_data[38934] <= r_data[38933];
                
                r_data[38935] <= r_data[38934];
                
                r_data[38936] <= r_data[38935];
                
                r_data[38937] <= r_data[38936];
                
                r_data[38938] <= r_data[38937];
                
                r_data[38939] <= r_data[38938];
                
                r_data[38940] <= r_data[38939];
                
                r_data[38941] <= r_data[38940];
                
                r_data[38942] <= r_data[38941];
                
                r_data[38943] <= r_data[38942];
                
                r_data[38944] <= r_data[38943];
                
                r_data[38945] <= r_data[38944];
                
                r_data[38946] <= r_data[38945];
                
                r_data[38947] <= r_data[38946];
                
                r_data[38948] <= r_data[38947];
                
                r_data[38949] <= r_data[38948];
                
                r_data[38950] <= r_data[38949];
                
                r_data[38951] <= r_data[38950];
                
                r_data[38952] <= r_data[38951];
                
                r_data[38953] <= r_data[38952];
                
                r_data[38954] <= r_data[38953];
                
                r_data[38955] <= r_data[38954];
                
                r_data[38956] <= r_data[38955];
                
                r_data[38957] <= r_data[38956];
                
                r_data[38958] <= r_data[38957];
                
                r_data[38959] <= r_data[38958];
                
                r_data[38960] <= r_data[38959];
                
                r_data[38961] <= r_data[38960];
                
                r_data[38962] <= r_data[38961];
                
                r_data[38963] <= r_data[38962];
                
                r_data[38964] <= r_data[38963];
                
                r_data[38965] <= r_data[38964];
                
                r_data[38966] <= r_data[38965];
                
                r_data[38967] <= r_data[38966];
                
                r_data[38968] <= r_data[38967];
                
                r_data[38969] <= r_data[38968];
                
                r_data[38970] <= r_data[38969];
                
                r_data[38971] <= r_data[38970];
                
                r_data[38972] <= r_data[38971];
                
                r_data[38973] <= r_data[38972];
                
                r_data[38974] <= r_data[38973];
                
                r_data[38975] <= r_data[38974];
                
                r_data[38976] <= r_data[38975];
                
                r_data[38977] <= r_data[38976];
                
                r_data[38978] <= r_data[38977];
                
                r_data[38979] <= r_data[38978];
                
                r_data[38980] <= r_data[38979];
                
                r_data[38981] <= r_data[38980];
                
                r_data[38982] <= r_data[38981];
                
                r_data[38983] <= r_data[38982];
                
                r_data[38984] <= r_data[38983];
                
                r_data[38985] <= r_data[38984];
                
                r_data[38986] <= r_data[38985];
                
                r_data[38987] <= r_data[38986];
                
                r_data[38988] <= r_data[38987];
                
                r_data[38989] <= r_data[38988];
                
                r_data[38990] <= r_data[38989];
                
                r_data[38991] <= r_data[38990];
                
                r_data[38992] <= r_data[38991];
                
                r_data[38993] <= r_data[38992];
                
                r_data[38994] <= r_data[38993];
                
                r_data[38995] <= r_data[38994];
                
                r_data[38996] <= r_data[38995];
                
                r_data[38997] <= r_data[38996];
                
                r_data[38998] <= r_data[38997];
                
                r_data[38999] <= r_data[38998];
                
                r_data[39000] <= r_data[38999];
                
                r_data[39001] <= r_data[39000];
                
                r_data[39002] <= r_data[39001];
                
                r_data[39003] <= r_data[39002];
                
                r_data[39004] <= r_data[39003];
                
                r_data[39005] <= r_data[39004];
                
                r_data[39006] <= r_data[39005];
                
                r_data[39007] <= r_data[39006];
                
                r_data[39008] <= r_data[39007];
                
                r_data[39009] <= r_data[39008];
                
                r_data[39010] <= r_data[39009];
                
                r_data[39011] <= r_data[39010];
                
                r_data[39012] <= r_data[39011];
                
                r_data[39013] <= r_data[39012];
                
                r_data[39014] <= r_data[39013];
                
                r_data[39015] <= r_data[39014];
                
                r_data[39016] <= r_data[39015];
                
                r_data[39017] <= r_data[39016];
                
                r_data[39018] <= r_data[39017];
                
                r_data[39019] <= r_data[39018];
                
                r_data[39020] <= r_data[39019];
                
                r_data[39021] <= r_data[39020];
                
                r_data[39022] <= r_data[39021];
                
                r_data[39023] <= r_data[39022];
                
                r_data[39024] <= r_data[39023];
                
                r_data[39025] <= r_data[39024];
                
                r_data[39026] <= r_data[39025];
                
                r_data[39027] <= r_data[39026];
                
                r_data[39028] <= r_data[39027];
                
                r_data[39029] <= r_data[39028];
                
                r_data[39030] <= r_data[39029];
                
                r_data[39031] <= r_data[39030];
                
                r_data[39032] <= r_data[39031];
                
                r_data[39033] <= r_data[39032];
                
                r_data[39034] <= r_data[39033];
                
                r_data[39035] <= r_data[39034];
                
                r_data[39036] <= r_data[39035];
                
                r_data[39037] <= r_data[39036];
                
                r_data[39038] <= r_data[39037];
                
                r_data[39039] <= r_data[39038];
                
                r_data[39040] <= r_data[39039];
                
                r_data[39041] <= r_data[39040];
                
                r_data[39042] <= r_data[39041];
                
                r_data[39043] <= r_data[39042];
                
                r_data[39044] <= r_data[39043];
                
                r_data[39045] <= r_data[39044];
                
                r_data[39046] <= r_data[39045];
                
                r_data[39047] <= r_data[39046];
                
                r_data[39048] <= r_data[39047];
                
                r_data[39049] <= r_data[39048];
                
                r_data[39050] <= r_data[39049];
                
                r_data[39051] <= r_data[39050];
                
                r_data[39052] <= r_data[39051];
                
                r_data[39053] <= r_data[39052];
                
                r_data[39054] <= r_data[39053];
                
                r_data[39055] <= r_data[39054];
                
                r_data[39056] <= r_data[39055];
                
                r_data[39057] <= r_data[39056];
                
                r_data[39058] <= r_data[39057];
                
                r_data[39059] <= r_data[39058];
                
                r_data[39060] <= r_data[39059];
                
                r_data[39061] <= r_data[39060];
                
                r_data[39062] <= r_data[39061];
                
                r_data[39063] <= r_data[39062];
                
                r_data[39064] <= r_data[39063];
                
                r_data[39065] <= r_data[39064];
                
                r_data[39066] <= r_data[39065];
                
                r_data[39067] <= r_data[39066];
                
                r_data[39068] <= r_data[39067];
                
                r_data[39069] <= r_data[39068];
                
                r_data[39070] <= r_data[39069];
                
                r_data[39071] <= r_data[39070];
                
                r_data[39072] <= r_data[39071];
                
                r_data[39073] <= r_data[39072];
                
                r_data[39074] <= r_data[39073];
                
                r_data[39075] <= r_data[39074];
                
                r_data[39076] <= r_data[39075];
                
                r_data[39077] <= r_data[39076];
                
                r_data[39078] <= r_data[39077];
                
                r_data[39079] <= r_data[39078];
                
                r_data[39080] <= r_data[39079];
                
                r_data[39081] <= r_data[39080];
                
                r_data[39082] <= r_data[39081];
                
                r_data[39083] <= r_data[39082];
                
                r_data[39084] <= r_data[39083];
                
                r_data[39085] <= r_data[39084];
                
                r_data[39086] <= r_data[39085];
                
                r_data[39087] <= r_data[39086];
                
                r_data[39088] <= r_data[39087];
                
                r_data[39089] <= r_data[39088];
                
                r_data[39090] <= r_data[39089];
                
                r_data[39091] <= r_data[39090];
                
                r_data[39092] <= r_data[39091];
                
                r_data[39093] <= r_data[39092];
                
                r_data[39094] <= r_data[39093];
                
                r_data[39095] <= r_data[39094];
                
                r_data[39096] <= r_data[39095];
                
                r_data[39097] <= r_data[39096];
                
                r_data[39098] <= r_data[39097];
                
                r_data[39099] <= r_data[39098];
                
                r_data[39100] <= r_data[39099];
                
                r_data[39101] <= r_data[39100];
                
                r_data[39102] <= r_data[39101];
                
                r_data[39103] <= r_data[39102];
                
                r_data[39104] <= r_data[39103];
                
                r_data[39105] <= r_data[39104];
                
                r_data[39106] <= r_data[39105];
                
                r_data[39107] <= r_data[39106];
                
                r_data[39108] <= r_data[39107];
                
                r_data[39109] <= r_data[39108];
                
                r_data[39110] <= r_data[39109];
                
                r_data[39111] <= r_data[39110];
                
                r_data[39112] <= r_data[39111];
                
                r_data[39113] <= r_data[39112];
                
                r_data[39114] <= r_data[39113];
                
                r_data[39115] <= r_data[39114];
                
                r_data[39116] <= r_data[39115];
                
                r_data[39117] <= r_data[39116];
                
                r_data[39118] <= r_data[39117];
                
                r_data[39119] <= r_data[39118];
                
                r_data[39120] <= r_data[39119];
                
                r_data[39121] <= r_data[39120];
                
                r_data[39122] <= r_data[39121];
                
                r_data[39123] <= r_data[39122];
                
                r_data[39124] <= r_data[39123];
                
                r_data[39125] <= r_data[39124];
                
                r_data[39126] <= r_data[39125];
                
                r_data[39127] <= r_data[39126];
                
                r_data[39128] <= r_data[39127];
                
                r_data[39129] <= r_data[39128];
                
                r_data[39130] <= r_data[39129];
                
                r_data[39131] <= r_data[39130];
                
                r_data[39132] <= r_data[39131];
                
                r_data[39133] <= r_data[39132];
                
                r_data[39134] <= r_data[39133];
                
                r_data[39135] <= r_data[39134];
                
                r_data[39136] <= r_data[39135];
                
                r_data[39137] <= r_data[39136];
                
                r_data[39138] <= r_data[39137];
                
                r_data[39139] <= r_data[39138];
                
                r_data[39140] <= r_data[39139];
                
                r_data[39141] <= r_data[39140];
                
                r_data[39142] <= r_data[39141];
                
                r_data[39143] <= r_data[39142];
                
                r_data[39144] <= r_data[39143];
                
                r_data[39145] <= r_data[39144];
                
                r_data[39146] <= r_data[39145];
                
                r_data[39147] <= r_data[39146];
                
                r_data[39148] <= r_data[39147];
                
                r_data[39149] <= r_data[39148];
                
                r_data[39150] <= r_data[39149];
                
                r_data[39151] <= r_data[39150];
                
                r_data[39152] <= r_data[39151];
                
                r_data[39153] <= r_data[39152];
                
                r_data[39154] <= r_data[39153];
                
                r_data[39155] <= r_data[39154];
                
                r_data[39156] <= r_data[39155];
                
                r_data[39157] <= r_data[39156];
                
                r_data[39158] <= r_data[39157];
                
                r_data[39159] <= r_data[39158];
                
                r_data[39160] <= r_data[39159];
                
                r_data[39161] <= r_data[39160];
                
                r_data[39162] <= r_data[39161];
                
                r_data[39163] <= r_data[39162];
                
                r_data[39164] <= r_data[39163];
                
                r_data[39165] <= r_data[39164];
                
                r_data[39166] <= r_data[39165];
                
                r_data[39167] <= r_data[39166];
                
                r_data[39168] <= r_data[39167];
                
                r_data[39169] <= r_data[39168];
                
                r_data[39170] <= r_data[39169];
                
                r_data[39171] <= r_data[39170];
                
                r_data[39172] <= r_data[39171];
                
                r_data[39173] <= r_data[39172];
                
                r_data[39174] <= r_data[39173];
                
                r_data[39175] <= r_data[39174];
                
                r_data[39176] <= r_data[39175];
                
                r_data[39177] <= r_data[39176];
                
                r_data[39178] <= r_data[39177];
                
                r_data[39179] <= r_data[39178];
                
                r_data[39180] <= r_data[39179];
                
                r_data[39181] <= r_data[39180];
                
                r_data[39182] <= r_data[39181];
                
                r_data[39183] <= r_data[39182];
                
                r_data[39184] <= r_data[39183];
                
                r_data[39185] <= r_data[39184];
                
                r_data[39186] <= r_data[39185];
                
                r_data[39187] <= r_data[39186];
                
                r_data[39188] <= r_data[39187];
                
                r_data[39189] <= r_data[39188];
                
                r_data[39190] <= r_data[39189];
                
                r_data[39191] <= r_data[39190];
                
                r_data[39192] <= r_data[39191];
                
                r_data[39193] <= r_data[39192];
                
                r_data[39194] <= r_data[39193];
                
                r_data[39195] <= r_data[39194];
                
                r_data[39196] <= r_data[39195];
                
                r_data[39197] <= r_data[39196];
                
                r_data[39198] <= r_data[39197];
                
                r_data[39199] <= r_data[39198];
                
                r_data[39200] <= r_data[39199];
                
                r_data[39201] <= r_data[39200];
                
                r_data[39202] <= r_data[39201];
                
                r_data[39203] <= r_data[39202];
                
                r_data[39204] <= r_data[39203];
                
                r_data[39205] <= r_data[39204];
                
                r_data[39206] <= r_data[39205];
                
                r_data[39207] <= r_data[39206];
                
                r_data[39208] <= r_data[39207];
                
                r_data[39209] <= r_data[39208];
                
                r_data[39210] <= r_data[39209];
                
                r_data[39211] <= r_data[39210];
                
                r_data[39212] <= r_data[39211];
                
                r_data[39213] <= r_data[39212];
                
                r_data[39214] <= r_data[39213];
                
                r_data[39215] <= r_data[39214];
                
                r_data[39216] <= r_data[39215];
                
                r_data[39217] <= r_data[39216];
                
                r_data[39218] <= r_data[39217];
                
                r_data[39219] <= r_data[39218];
                
                r_data[39220] <= r_data[39219];
                
                r_data[39221] <= r_data[39220];
                
                r_data[39222] <= r_data[39221];
                
                r_data[39223] <= r_data[39222];
                
                r_data[39224] <= r_data[39223];
                
                r_data[39225] <= r_data[39224];
                
                r_data[39226] <= r_data[39225];
                
                r_data[39227] <= r_data[39226];
                
                r_data[39228] <= r_data[39227];
                
                r_data[39229] <= r_data[39228];
                
                r_data[39230] <= r_data[39229];
                
                r_data[39231] <= r_data[39230];
                
                r_data[39232] <= r_data[39231];
                
                r_data[39233] <= r_data[39232];
                
                r_data[39234] <= r_data[39233];
                
                r_data[39235] <= r_data[39234];
                
                r_data[39236] <= r_data[39235];
                
                r_data[39237] <= r_data[39236];
                
                r_data[39238] <= r_data[39237];
                
                r_data[39239] <= r_data[39238];
                
                r_data[39240] <= r_data[39239];
                
                r_data[39241] <= r_data[39240];
                
                r_data[39242] <= r_data[39241];
                
                r_data[39243] <= r_data[39242];
                
                r_data[39244] <= r_data[39243];
                
                r_data[39245] <= r_data[39244];
                
                r_data[39246] <= r_data[39245];
                
                r_data[39247] <= r_data[39246];
                
                r_data[39248] <= r_data[39247];
                
                r_data[39249] <= r_data[39248];
                
                r_data[39250] <= r_data[39249];
                
                r_data[39251] <= r_data[39250];
                
                r_data[39252] <= r_data[39251];
                
                r_data[39253] <= r_data[39252];
                
                r_data[39254] <= r_data[39253];
                
                r_data[39255] <= r_data[39254];
                
                r_data[39256] <= r_data[39255];
                
                r_data[39257] <= r_data[39256];
                
                r_data[39258] <= r_data[39257];
                
                r_data[39259] <= r_data[39258];
                
                r_data[39260] <= r_data[39259];
                
                r_data[39261] <= r_data[39260];
                
                r_data[39262] <= r_data[39261];
                
                r_data[39263] <= r_data[39262];
                
                r_data[39264] <= r_data[39263];
                
                r_data[39265] <= r_data[39264];
                
                r_data[39266] <= r_data[39265];
                
                r_data[39267] <= r_data[39266];
                
                r_data[39268] <= r_data[39267];
                
                r_data[39269] <= r_data[39268];
                
                r_data[39270] <= r_data[39269];
                
                r_data[39271] <= r_data[39270];
                
                r_data[39272] <= r_data[39271];
                
                r_data[39273] <= r_data[39272];
                
                r_data[39274] <= r_data[39273];
                
                r_data[39275] <= r_data[39274];
                
                r_data[39276] <= r_data[39275];
                
                r_data[39277] <= r_data[39276];
                
                r_data[39278] <= r_data[39277];
                
                r_data[39279] <= r_data[39278];
                
                r_data[39280] <= r_data[39279];
                
                r_data[39281] <= r_data[39280];
                
                r_data[39282] <= r_data[39281];
                
                r_data[39283] <= r_data[39282];
                
                r_data[39284] <= r_data[39283];
                
                r_data[39285] <= r_data[39284];
                
                r_data[39286] <= r_data[39285];
                
                r_data[39287] <= r_data[39286];
                
                r_data[39288] <= r_data[39287];
                
                r_data[39289] <= r_data[39288];
                
                r_data[39290] <= r_data[39289];
                
                r_data[39291] <= r_data[39290];
                
                r_data[39292] <= r_data[39291];
                
                r_data[39293] <= r_data[39292];
                
                r_data[39294] <= r_data[39293];
                
                r_data[39295] <= r_data[39294];
                
                r_data[39296] <= r_data[39295];
                
                r_data[39297] <= r_data[39296];
                
                r_data[39298] <= r_data[39297];
                
                r_data[39299] <= r_data[39298];
                
                r_data[39300] <= r_data[39299];
                
                r_data[39301] <= r_data[39300];
                
                r_data[39302] <= r_data[39301];
                
                r_data[39303] <= r_data[39302];
                
                r_data[39304] <= r_data[39303];
                
                r_data[39305] <= r_data[39304];
                
                r_data[39306] <= r_data[39305];
                
                r_data[39307] <= r_data[39306];
                
                r_data[39308] <= r_data[39307];
                
                r_data[39309] <= r_data[39308];
                
                r_data[39310] <= r_data[39309];
                
                r_data[39311] <= r_data[39310];
                
                r_data[39312] <= r_data[39311];
                
                r_data[39313] <= r_data[39312];
                
                r_data[39314] <= r_data[39313];
                
                r_data[39315] <= r_data[39314];
                
                r_data[39316] <= r_data[39315];
                
                r_data[39317] <= r_data[39316];
                
                r_data[39318] <= r_data[39317];
                
                r_data[39319] <= r_data[39318];
                
                r_data[39320] <= r_data[39319];
                
                r_data[39321] <= r_data[39320];
                
                r_data[39322] <= r_data[39321];
                
                r_data[39323] <= r_data[39322];
                
                r_data[39324] <= r_data[39323];
                
                r_data[39325] <= r_data[39324];
                
                r_data[39326] <= r_data[39325];
                
                r_data[39327] <= r_data[39326];
                
                r_data[39328] <= r_data[39327];
                
                r_data[39329] <= r_data[39328];
                
                r_data[39330] <= r_data[39329];
                
                r_data[39331] <= r_data[39330];
                
                r_data[39332] <= r_data[39331];
                
                r_data[39333] <= r_data[39332];
                
                r_data[39334] <= r_data[39333];
                
                r_data[39335] <= r_data[39334];
                
                r_data[39336] <= r_data[39335];
                
                r_data[39337] <= r_data[39336];
                
                r_data[39338] <= r_data[39337];
                
                r_data[39339] <= r_data[39338];
                
                r_data[39340] <= r_data[39339];
                
                r_data[39341] <= r_data[39340];
                
                r_data[39342] <= r_data[39341];
                
                r_data[39343] <= r_data[39342];
                
                r_data[39344] <= r_data[39343];
                
                r_data[39345] <= r_data[39344];
                
                r_data[39346] <= r_data[39345];
                
                r_data[39347] <= r_data[39346];
                
                r_data[39348] <= r_data[39347];
                
                r_data[39349] <= r_data[39348];
                
                r_data[39350] <= r_data[39349];
                
                r_data[39351] <= r_data[39350];
                
                r_data[39352] <= r_data[39351];
                
                r_data[39353] <= r_data[39352];
                
                r_data[39354] <= r_data[39353];
                
                r_data[39355] <= r_data[39354];
                
                r_data[39356] <= r_data[39355];
                
                r_data[39357] <= r_data[39356];
                
                r_data[39358] <= r_data[39357];
                
                r_data[39359] <= r_data[39358];
                
                r_data[39360] <= r_data[39359];
                
                r_data[39361] <= r_data[39360];
                
                r_data[39362] <= r_data[39361];
                
                r_data[39363] <= r_data[39362];
                
                r_data[39364] <= r_data[39363];
                
                r_data[39365] <= r_data[39364];
                
                r_data[39366] <= r_data[39365];
                
                r_data[39367] <= r_data[39366];
                
                r_data[39368] <= r_data[39367];
                
                r_data[39369] <= r_data[39368];
                
                r_data[39370] <= r_data[39369];
                
                r_data[39371] <= r_data[39370];
                
                r_data[39372] <= r_data[39371];
                
                r_data[39373] <= r_data[39372];
                
                r_data[39374] <= r_data[39373];
                
                r_data[39375] <= r_data[39374];
                
                r_data[39376] <= r_data[39375];
                
                r_data[39377] <= r_data[39376];
                
                r_data[39378] <= r_data[39377];
                
                r_data[39379] <= r_data[39378];
                
                r_data[39380] <= r_data[39379];
                
                r_data[39381] <= r_data[39380];
                
                r_data[39382] <= r_data[39381];
                
                r_data[39383] <= r_data[39382];
                
                r_data[39384] <= r_data[39383];
                
                r_data[39385] <= r_data[39384];
                
                r_data[39386] <= r_data[39385];
                
                r_data[39387] <= r_data[39386];
                
                r_data[39388] <= r_data[39387];
                
                r_data[39389] <= r_data[39388];
                
                r_data[39390] <= r_data[39389];
                
                r_data[39391] <= r_data[39390];
                
                r_data[39392] <= r_data[39391];
                
                r_data[39393] <= r_data[39392];
                
                r_data[39394] <= r_data[39393];
                
                r_data[39395] <= r_data[39394];
                
                r_data[39396] <= r_data[39395];
                
                r_data[39397] <= r_data[39396];
                
                r_data[39398] <= r_data[39397];
                
                r_data[39399] <= r_data[39398];
                
                r_data[39400] <= r_data[39399];
                
                r_data[39401] <= r_data[39400];
                
                r_data[39402] <= r_data[39401];
                
                r_data[39403] <= r_data[39402];
                
                r_data[39404] <= r_data[39403];
                
                r_data[39405] <= r_data[39404];
                
                r_data[39406] <= r_data[39405];
                
                r_data[39407] <= r_data[39406];
                
                r_data[39408] <= r_data[39407];
                
                r_data[39409] <= r_data[39408];
                
                r_data[39410] <= r_data[39409];
                
                r_data[39411] <= r_data[39410];
                
                r_data[39412] <= r_data[39411];
                
                r_data[39413] <= r_data[39412];
                
                r_data[39414] <= r_data[39413];
                
                r_data[39415] <= r_data[39414];
                
                r_data[39416] <= r_data[39415];
                
                r_data[39417] <= r_data[39416];
                
                r_data[39418] <= r_data[39417];
                
                r_data[39419] <= r_data[39418];
                
                r_data[39420] <= r_data[39419];
                
                r_data[39421] <= r_data[39420];
                
                r_data[39422] <= r_data[39421];
                
                r_data[39423] <= r_data[39422];
                
                r_data[39424] <= r_data[39423];
                
                r_data[39425] <= r_data[39424];
                
                r_data[39426] <= r_data[39425];
                
                r_data[39427] <= r_data[39426];
                
                r_data[39428] <= r_data[39427];
                
                r_data[39429] <= r_data[39428];
                
                r_data[39430] <= r_data[39429];
                
                r_data[39431] <= r_data[39430];
                
                r_data[39432] <= r_data[39431];
                
                r_data[39433] <= r_data[39432];
                
                r_data[39434] <= r_data[39433];
                
                r_data[39435] <= r_data[39434];
                
                r_data[39436] <= r_data[39435];
                
                r_data[39437] <= r_data[39436];
                
                r_data[39438] <= r_data[39437];
                
                r_data[39439] <= r_data[39438];
                
                r_data[39440] <= r_data[39439];
                
                r_data[39441] <= r_data[39440];
                
                r_data[39442] <= r_data[39441];
                
                r_data[39443] <= r_data[39442];
                
                r_data[39444] <= r_data[39443];
                
                r_data[39445] <= r_data[39444];
                
                r_data[39446] <= r_data[39445];
                
                r_data[39447] <= r_data[39446];
                
                r_data[39448] <= r_data[39447];
                
                r_data[39449] <= r_data[39448];
                
                r_data[39450] <= r_data[39449];
                
                r_data[39451] <= r_data[39450];
                
                r_data[39452] <= r_data[39451];
                
                r_data[39453] <= r_data[39452];
                
                r_data[39454] <= r_data[39453];
                
                r_data[39455] <= r_data[39454];
                
                r_data[39456] <= r_data[39455];
                
                r_data[39457] <= r_data[39456];
                
                r_data[39458] <= r_data[39457];
                
                r_data[39459] <= r_data[39458];
                
                r_data[39460] <= r_data[39459];
                
                r_data[39461] <= r_data[39460];
                
                r_data[39462] <= r_data[39461];
                
                r_data[39463] <= r_data[39462];
                
                r_data[39464] <= r_data[39463];
                
                r_data[39465] <= r_data[39464];
                
                r_data[39466] <= r_data[39465];
                
                r_data[39467] <= r_data[39466];
                
                r_data[39468] <= r_data[39467];
                
                r_data[39469] <= r_data[39468];
                
                r_data[39470] <= r_data[39469];
                
                r_data[39471] <= r_data[39470];
                
                r_data[39472] <= r_data[39471];
                
                r_data[39473] <= r_data[39472];
                
                r_data[39474] <= r_data[39473];
                
                r_data[39475] <= r_data[39474];
                
                r_data[39476] <= r_data[39475];
                
                r_data[39477] <= r_data[39476];
                
                r_data[39478] <= r_data[39477];
                
                r_data[39479] <= r_data[39478];
                
                r_data[39480] <= r_data[39479];
                
                r_data[39481] <= r_data[39480];
                
                r_data[39482] <= r_data[39481];
                
                r_data[39483] <= r_data[39482];
                
                r_data[39484] <= r_data[39483];
                
                r_data[39485] <= r_data[39484];
                
                r_data[39486] <= r_data[39485];
                
                r_data[39487] <= r_data[39486];
                
                r_data[39488] <= r_data[39487];
                
                r_data[39489] <= r_data[39488];
                
                r_data[39490] <= r_data[39489];
                
                r_data[39491] <= r_data[39490];
                
                r_data[39492] <= r_data[39491];
                
                r_data[39493] <= r_data[39492];
                
                r_data[39494] <= r_data[39493];
                
                r_data[39495] <= r_data[39494];
                
                r_data[39496] <= r_data[39495];
                
                r_data[39497] <= r_data[39496];
                
                r_data[39498] <= r_data[39497];
                
                r_data[39499] <= r_data[39498];
                
                r_data[39500] <= r_data[39499];
                
                r_data[39501] <= r_data[39500];
                
                r_data[39502] <= r_data[39501];
                
                r_data[39503] <= r_data[39502];
                
                r_data[39504] <= r_data[39503];
                
                r_data[39505] <= r_data[39504];
                
                r_data[39506] <= r_data[39505];
                
                r_data[39507] <= r_data[39506];
                
                r_data[39508] <= r_data[39507];
                
                r_data[39509] <= r_data[39508];
                
                r_data[39510] <= r_data[39509];
                
                r_data[39511] <= r_data[39510];
                
                r_data[39512] <= r_data[39511];
                
                r_data[39513] <= r_data[39512];
                
                r_data[39514] <= r_data[39513];
                
                r_data[39515] <= r_data[39514];
                
                r_data[39516] <= r_data[39515];
                
                r_data[39517] <= r_data[39516];
                
                r_data[39518] <= r_data[39517];
                
                r_data[39519] <= r_data[39518];
                
                r_data[39520] <= r_data[39519];
                
                r_data[39521] <= r_data[39520];
                
                r_data[39522] <= r_data[39521];
                
                r_data[39523] <= r_data[39522];
                
                r_data[39524] <= r_data[39523];
                
                r_data[39525] <= r_data[39524];
                
                r_data[39526] <= r_data[39525];
                
                r_data[39527] <= r_data[39526];
                
                r_data[39528] <= r_data[39527];
                
                r_data[39529] <= r_data[39528];
                
                r_data[39530] <= r_data[39529];
                
                r_data[39531] <= r_data[39530];
                
                r_data[39532] <= r_data[39531];
                
                r_data[39533] <= r_data[39532];
                
                r_data[39534] <= r_data[39533];
                
                r_data[39535] <= r_data[39534];
                
                r_data[39536] <= r_data[39535];
                
                r_data[39537] <= r_data[39536];
                
                r_data[39538] <= r_data[39537];
                
                r_data[39539] <= r_data[39538];
                
                r_data[39540] <= r_data[39539];
                
                r_data[39541] <= r_data[39540];
                
                r_data[39542] <= r_data[39541];
                
                r_data[39543] <= r_data[39542];
                
                r_data[39544] <= r_data[39543];
                
                r_data[39545] <= r_data[39544];
                
                r_data[39546] <= r_data[39545];
                
                r_data[39547] <= r_data[39546];
                
                r_data[39548] <= r_data[39547];
                
                r_data[39549] <= r_data[39548];
                
                r_data[39550] <= r_data[39549];
                
                r_data[39551] <= r_data[39550];
                
                r_data[39552] <= r_data[39551];
                
                r_data[39553] <= r_data[39552];
                
                r_data[39554] <= r_data[39553];
                
                r_data[39555] <= r_data[39554];
                
                r_data[39556] <= r_data[39555];
                
                r_data[39557] <= r_data[39556];
                
                r_data[39558] <= r_data[39557];
                
                r_data[39559] <= r_data[39558];
                
                r_data[39560] <= r_data[39559];
                
                r_data[39561] <= r_data[39560];
                
                r_data[39562] <= r_data[39561];
                
                r_data[39563] <= r_data[39562];
                
                r_data[39564] <= r_data[39563];
                
                r_data[39565] <= r_data[39564];
                
                r_data[39566] <= r_data[39565];
                
                r_data[39567] <= r_data[39566];
                
                r_data[39568] <= r_data[39567];
                
                r_data[39569] <= r_data[39568];
                
                r_data[39570] <= r_data[39569];
                
                r_data[39571] <= r_data[39570];
                
                r_data[39572] <= r_data[39571];
                
                r_data[39573] <= r_data[39572];
                
                r_data[39574] <= r_data[39573];
                
                r_data[39575] <= r_data[39574];
                
                r_data[39576] <= r_data[39575];
                
                r_data[39577] <= r_data[39576];
                
                r_data[39578] <= r_data[39577];
                
                r_data[39579] <= r_data[39578];
                
                r_data[39580] <= r_data[39579];
                
                r_data[39581] <= r_data[39580];
                
                r_data[39582] <= r_data[39581];
                
                r_data[39583] <= r_data[39582];
                
                r_data[39584] <= r_data[39583];
                
                r_data[39585] <= r_data[39584];
                
                r_data[39586] <= r_data[39585];
                
                r_data[39587] <= r_data[39586];
                
                r_data[39588] <= r_data[39587];
                
                r_data[39589] <= r_data[39588];
                
                r_data[39590] <= r_data[39589];
                
                r_data[39591] <= r_data[39590];
                
                r_data[39592] <= r_data[39591];
                
                r_data[39593] <= r_data[39592];
                
                r_data[39594] <= r_data[39593];
                
                r_data[39595] <= r_data[39594];
                
                r_data[39596] <= r_data[39595];
                
                r_data[39597] <= r_data[39596];
                
                r_data[39598] <= r_data[39597];
                
                r_data[39599] <= r_data[39598];
                
                r_data[39600] <= r_data[39599];
                
                r_data[39601] <= r_data[39600];
                
                r_data[39602] <= r_data[39601];
                
                r_data[39603] <= r_data[39602];
                
                r_data[39604] <= r_data[39603];
                
                r_data[39605] <= r_data[39604];
                
                r_data[39606] <= r_data[39605];
                
                r_data[39607] <= r_data[39606];
                
                r_data[39608] <= r_data[39607];
                
                r_data[39609] <= r_data[39608];
                
                r_data[39610] <= r_data[39609];
                
                r_data[39611] <= r_data[39610];
                
                r_data[39612] <= r_data[39611];
                
                r_data[39613] <= r_data[39612];
                
                r_data[39614] <= r_data[39613];
                
                r_data[39615] <= r_data[39614];
                
                r_data[39616] <= r_data[39615];
                
                r_data[39617] <= r_data[39616];
                
                r_data[39618] <= r_data[39617];
                
                r_data[39619] <= r_data[39618];
                
                r_data[39620] <= r_data[39619];
                
                r_data[39621] <= r_data[39620];
                
                r_data[39622] <= r_data[39621];
                
                r_data[39623] <= r_data[39622];
                
                r_data[39624] <= r_data[39623];
                
                r_data[39625] <= r_data[39624];
                
                r_data[39626] <= r_data[39625];
                
                r_data[39627] <= r_data[39626];
                
                r_data[39628] <= r_data[39627];
                
                r_data[39629] <= r_data[39628];
                
                r_data[39630] <= r_data[39629];
                
                r_data[39631] <= r_data[39630];
                
                r_data[39632] <= r_data[39631];
                
                r_data[39633] <= r_data[39632];
                
                r_data[39634] <= r_data[39633];
                
                r_data[39635] <= r_data[39634];
                
                r_data[39636] <= r_data[39635];
                
                r_data[39637] <= r_data[39636];
                
                r_data[39638] <= r_data[39637];
                
                r_data[39639] <= r_data[39638];
                
                r_data[39640] <= r_data[39639];
                
                r_data[39641] <= r_data[39640];
                
                r_data[39642] <= r_data[39641];
                
                r_data[39643] <= r_data[39642];
                
                r_data[39644] <= r_data[39643];
                
                r_data[39645] <= r_data[39644];
                
                r_data[39646] <= r_data[39645];
                
                r_data[39647] <= r_data[39646];
                
                r_data[39648] <= r_data[39647];
                
                r_data[39649] <= r_data[39648];
                
                r_data[39650] <= r_data[39649];
                
                r_data[39651] <= r_data[39650];
                
                r_data[39652] <= r_data[39651];
                
                r_data[39653] <= r_data[39652];
                
                r_data[39654] <= r_data[39653];
                
                r_data[39655] <= r_data[39654];
                
                r_data[39656] <= r_data[39655];
                
                r_data[39657] <= r_data[39656];
                
                r_data[39658] <= r_data[39657];
                
                r_data[39659] <= r_data[39658];
                
                r_data[39660] <= r_data[39659];
                
                r_data[39661] <= r_data[39660];
                
                r_data[39662] <= r_data[39661];
                
                r_data[39663] <= r_data[39662];
                
                r_data[39664] <= r_data[39663];
                
                r_data[39665] <= r_data[39664];
                
                r_data[39666] <= r_data[39665];
                
                r_data[39667] <= r_data[39666];
                
                r_data[39668] <= r_data[39667];
                
                r_data[39669] <= r_data[39668];
                
                r_data[39670] <= r_data[39669];
                
                r_data[39671] <= r_data[39670];
                
                r_data[39672] <= r_data[39671];
                
                r_data[39673] <= r_data[39672];
                
                r_data[39674] <= r_data[39673];
                
                r_data[39675] <= r_data[39674];
                
                r_data[39676] <= r_data[39675];
                
                r_data[39677] <= r_data[39676];
                
                r_data[39678] <= r_data[39677];
                
                r_data[39679] <= r_data[39678];
                
                r_data[39680] <= r_data[39679];
                
                r_data[39681] <= r_data[39680];
                
                r_data[39682] <= r_data[39681];
                
                r_data[39683] <= r_data[39682];
                
                r_data[39684] <= r_data[39683];
                
                r_data[39685] <= r_data[39684];
                
                r_data[39686] <= r_data[39685];
                
                r_data[39687] <= r_data[39686];
                
                r_data[39688] <= r_data[39687];
                
                r_data[39689] <= r_data[39688];
                
                r_data[39690] <= r_data[39689];
                
                r_data[39691] <= r_data[39690];
                
                r_data[39692] <= r_data[39691];
                
                r_data[39693] <= r_data[39692];
                
                r_data[39694] <= r_data[39693];
                
                r_data[39695] <= r_data[39694];
                
                r_data[39696] <= r_data[39695];
                
                r_data[39697] <= r_data[39696];
                
                r_data[39698] <= r_data[39697];
                
                r_data[39699] <= r_data[39698];
                
                r_data[39700] <= r_data[39699];
                
                r_data[39701] <= r_data[39700];
                
                r_data[39702] <= r_data[39701];
                
                r_data[39703] <= r_data[39702];
                
                r_data[39704] <= r_data[39703];
                
                r_data[39705] <= r_data[39704];
                
                r_data[39706] <= r_data[39705];
                
                r_data[39707] <= r_data[39706];
                
                r_data[39708] <= r_data[39707];
                
                r_data[39709] <= r_data[39708];
                
                r_data[39710] <= r_data[39709];
                
                r_data[39711] <= r_data[39710];
                
                r_data[39712] <= r_data[39711];
                
                r_data[39713] <= r_data[39712];
                
                r_data[39714] <= r_data[39713];
                
                r_data[39715] <= r_data[39714];
                
                r_data[39716] <= r_data[39715];
                
                r_data[39717] <= r_data[39716];
                
                r_data[39718] <= r_data[39717];
                
                r_data[39719] <= r_data[39718];
                
                r_data[39720] <= r_data[39719];
                
                r_data[39721] <= r_data[39720];
                
                r_data[39722] <= r_data[39721];
                
                r_data[39723] <= r_data[39722];
                
                r_data[39724] <= r_data[39723];
                
                r_data[39725] <= r_data[39724];
                
                r_data[39726] <= r_data[39725];
                
                r_data[39727] <= r_data[39726];
                
                r_data[39728] <= r_data[39727];
                
                r_data[39729] <= r_data[39728];
                
                r_data[39730] <= r_data[39729];
                
                r_data[39731] <= r_data[39730];
                
                r_data[39732] <= r_data[39731];
                
                r_data[39733] <= r_data[39732];
                
                r_data[39734] <= r_data[39733];
                
                r_data[39735] <= r_data[39734];
                
                r_data[39736] <= r_data[39735];
                
                r_data[39737] <= r_data[39736];
                
                r_data[39738] <= r_data[39737];
                
                r_data[39739] <= r_data[39738];
                
                r_data[39740] <= r_data[39739];
                
                r_data[39741] <= r_data[39740];
                
                r_data[39742] <= r_data[39741];
                
                r_data[39743] <= r_data[39742];
                
                r_data[39744] <= r_data[39743];
                
                r_data[39745] <= r_data[39744];
                
                r_data[39746] <= r_data[39745];
                
                r_data[39747] <= r_data[39746];
                
                r_data[39748] <= r_data[39747];
                
                r_data[39749] <= r_data[39748];
                
                r_data[39750] <= r_data[39749];
                
                r_data[39751] <= r_data[39750];
                
                r_data[39752] <= r_data[39751];
                
                r_data[39753] <= r_data[39752];
                
                r_data[39754] <= r_data[39753];
                
                r_data[39755] <= r_data[39754];
                
                r_data[39756] <= r_data[39755];
                
                r_data[39757] <= r_data[39756];
                
                r_data[39758] <= r_data[39757];
                
                r_data[39759] <= r_data[39758];
                
                r_data[39760] <= r_data[39759];
                
                r_data[39761] <= r_data[39760];
                
                r_data[39762] <= r_data[39761];
                
                r_data[39763] <= r_data[39762];
                
                r_data[39764] <= r_data[39763];
                
                r_data[39765] <= r_data[39764];
                
                r_data[39766] <= r_data[39765];
                
                r_data[39767] <= r_data[39766];
                
                r_data[39768] <= r_data[39767];
                
                r_data[39769] <= r_data[39768];
                
                r_data[39770] <= r_data[39769];
                
                r_data[39771] <= r_data[39770];
                
                r_data[39772] <= r_data[39771];
                
                r_data[39773] <= r_data[39772];
                
                r_data[39774] <= r_data[39773];
                
                r_data[39775] <= r_data[39774];
                
                r_data[39776] <= r_data[39775];
                
                r_data[39777] <= r_data[39776];
                
                r_data[39778] <= r_data[39777];
                
                r_data[39779] <= r_data[39778];
                
                r_data[39780] <= r_data[39779];
                
                r_data[39781] <= r_data[39780];
                
                r_data[39782] <= r_data[39781];
                
                r_data[39783] <= r_data[39782];
                
                r_data[39784] <= r_data[39783];
                
                r_data[39785] <= r_data[39784];
                
                r_data[39786] <= r_data[39785];
                
                r_data[39787] <= r_data[39786];
                
                r_data[39788] <= r_data[39787];
                
                r_data[39789] <= r_data[39788];
                
                r_data[39790] <= r_data[39789];
                
                r_data[39791] <= r_data[39790];
                
                r_data[39792] <= r_data[39791];
                
                r_data[39793] <= r_data[39792];
                
                r_data[39794] <= r_data[39793];
                
                r_data[39795] <= r_data[39794];
                
                r_data[39796] <= r_data[39795];
                
                r_data[39797] <= r_data[39796];
                
                r_data[39798] <= r_data[39797];
                
                r_data[39799] <= r_data[39798];
                
                r_data[39800] <= r_data[39799];
                
                r_data[39801] <= r_data[39800];
                
                r_data[39802] <= r_data[39801];
                
                r_data[39803] <= r_data[39802];
                
                r_data[39804] <= r_data[39803];
                
                r_data[39805] <= r_data[39804];
                
                r_data[39806] <= r_data[39805];
                
                r_data[39807] <= r_data[39806];
                
                r_data[39808] <= r_data[39807];
                
                r_data[39809] <= r_data[39808];
                
                r_data[39810] <= r_data[39809];
                
                r_data[39811] <= r_data[39810];
                
                r_data[39812] <= r_data[39811];
                
                r_data[39813] <= r_data[39812];
                
                r_data[39814] <= r_data[39813];
                
                r_data[39815] <= r_data[39814];
                
                r_data[39816] <= r_data[39815];
                
                r_data[39817] <= r_data[39816];
                
                r_data[39818] <= r_data[39817];
                
                r_data[39819] <= r_data[39818];
                
                r_data[39820] <= r_data[39819];
                
                r_data[39821] <= r_data[39820];
                
                r_data[39822] <= r_data[39821];
                
                r_data[39823] <= r_data[39822];
                
                r_data[39824] <= r_data[39823];
                
                r_data[39825] <= r_data[39824];
                
                r_data[39826] <= r_data[39825];
                
                r_data[39827] <= r_data[39826];
                
                r_data[39828] <= r_data[39827];
                
                r_data[39829] <= r_data[39828];
                
                r_data[39830] <= r_data[39829];
                
                r_data[39831] <= r_data[39830];
                
                r_data[39832] <= r_data[39831];
                
                r_data[39833] <= r_data[39832];
                
                r_data[39834] <= r_data[39833];
                
                r_data[39835] <= r_data[39834];
                
                r_data[39836] <= r_data[39835];
                
                r_data[39837] <= r_data[39836];
                
                r_data[39838] <= r_data[39837];
                
                r_data[39839] <= r_data[39838];
                
                r_data[39840] <= r_data[39839];
                
                r_data[39841] <= r_data[39840];
                
                r_data[39842] <= r_data[39841];
                
                r_data[39843] <= r_data[39842];
                
                r_data[39844] <= r_data[39843];
                
                r_data[39845] <= r_data[39844];
                
                r_data[39846] <= r_data[39845];
                
                r_data[39847] <= r_data[39846];
                
                r_data[39848] <= r_data[39847];
                
                r_data[39849] <= r_data[39848];
                
                r_data[39850] <= r_data[39849];
                
                r_data[39851] <= r_data[39850];
                
                r_data[39852] <= r_data[39851];
                
                r_data[39853] <= r_data[39852];
                
                r_data[39854] <= r_data[39853];
                
                r_data[39855] <= r_data[39854];
                
                r_data[39856] <= r_data[39855];
                
                r_data[39857] <= r_data[39856];
                
                r_data[39858] <= r_data[39857];
                
                r_data[39859] <= r_data[39858];
                
                r_data[39860] <= r_data[39859];
                
                r_data[39861] <= r_data[39860];
                
                r_data[39862] <= r_data[39861];
                
                r_data[39863] <= r_data[39862];
                
                r_data[39864] <= r_data[39863];
                
                r_data[39865] <= r_data[39864];
                
                r_data[39866] <= r_data[39865];
                
                r_data[39867] <= r_data[39866];
                
                r_data[39868] <= r_data[39867];
                
                r_data[39869] <= r_data[39868];
                
                r_data[39870] <= r_data[39869];
                
                r_data[39871] <= r_data[39870];
                
                r_data[39872] <= r_data[39871];
                
                r_data[39873] <= r_data[39872];
                
                r_data[39874] <= r_data[39873];
                
                r_data[39875] <= r_data[39874];
                
                r_data[39876] <= r_data[39875];
                
                r_data[39877] <= r_data[39876];
                
                r_data[39878] <= r_data[39877];
                
                r_data[39879] <= r_data[39878];
                
                r_data[39880] <= r_data[39879];
                
                r_data[39881] <= r_data[39880];
                
                r_data[39882] <= r_data[39881];
                
                r_data[39883] <= r_data[39882];
                
                r_data[39884] <= r_data[39883];
                
                r_data[39885] <= r_data[39884];
                
                r_data[39886] <= r_data[39885];
                
                r_data[39887] <= r_data[39886];
                
                r_data[39888] <= r_data[39887];
                
                r_data[39889] <= r_data[39888];
                
                r_data[39890] <= r_data[39889];
                
                r_data[39891] <= r_data[39890];
                
                r_data[39892] <= r_data[39891];
                
                r_data[39893] <= r_data[39892];
                
                r_data[39894] <= r_data[39893];
                
                r_data[39895] <= r_data[39894];
                
                r_data[39896] <= r_data[39895];
                
                r_data[39897] <= r_data[39896];
                
                r_data[39898] <= r_data[39897];
                
                r_data[39899] <= r_data[39898];
                
                r_data[39900] <= r_data[39899];
                
                r_data[39901] <= r_data[39900];
                
                r_data[39902] <= r_data[39901];
                
                r_data[39903] <= r_data[39902];
                
                r_data[39904] <= r_data[39903];
                
                r_data[39905] <= r_data[39904];
                
                r_data[39906] <= r_data[39905];
                
                r_data[39907] <= r_data[39906];
                
                r_data[39908] <= r_data[39907];
                
                r_data[39909] <= r_data[39908];
                
                r_data[39910] <= r_data[39909];
                
                r_data[39911] <= r_data[39910];
                
                r_data[39912] <= r_data[39911];
                
                r_data[39913] <= r_data[39912];
                
                r_data[39914] <= r_data[39913];
                
                r_data[39915] <= r_data[39914];
                
                r_data[39916] <= r_data[39915];
                
                r_data[39917] <= r_data[39916];
                
                r_data[39918] <= r_data[39917];
                
                r_data[39919] <= r_data[39918];
                
                r_data[39920] <= r_data[39919];
                
                r_data[39921] <= r_data[39920];
                
                r_data[39922] <= r_data[39921];
                
                r_data[39923] <= r_data[39922];
                
                r_data[39924] <= r_data[39923];
                
                r_data[39925] <= r_data[39924];
                
                r_data[39926] <= r_data[39925];
                
                r_data[39927] <= r_data[39926];
                
                r_data[39928] <= r_data[39927];
                
                r_data[39929] <= r_data[39928];
                
                r_data[39930] <= r_data[39929];
                
                r_data[39931] <= r_data[39930];
                
                r_data[39932] <= r_data[39931];
                
                r_data[39933] <= r_data[39932];
                
                r_data[39934] <= r_data[39933];
                
                r_data[39935] <= r_data[39934];
                
                r_data[39936] <= r_data[39935];
                
                r_data[39937] <= r_data[39936];
                
                r_data[39938] <= r_data[39937];
                
                r_data[39939] <= r_data[39938];
                
                r_data[39940] <= r_data[39939];
                
                r_data[39941] <= r_data[39940];
                
                r_data[39942] <= r_data[39941];
                
                r_data[39943] <= r_data[39942];
                
                r_data[39944] <= r_data[39943];
                
                r_data[39945] <= r_data[39944];
                
                r_data[39946] <= r_data[39945];
                
                r_data[39947] <= r_data[39946];
                
                r_data[39948] <= r_data[39947];
                
                r_data[39949] <= r_data[39948];
                
                r_data[39950] <= r_data[39949];
                
                r_data[39951] <= r_data[39950];
                
                r_data[39952] <= r_data[39951];
                
                r_data[39953] <= r_data[39952];
                
                r_data[39954] <= r_data[39953];
                
                r_data[39955] <= r_data[39954];
                
                r_data[39956] <= r_data[39955];
                
                r_data[39957] <= r_data[39956];
                
                r_data[39958] <= r_data[39957];
                
                r_data[39959] <= r_data[39958];
                
                r_data[39960] <= r_data[39959];
                
                r_data[39961] <= r_data[39960];
                
                r_data[39962] <= r_data[39961];
                
                r_data[39963] <= r_data[39962];
                
                r_data[39964] <= r_data[39963];
                
                r_data[39965] <= r_data[39964];
                
                r_data[39966] <= r_data[39965];
                
                r_data[39967] <= r_data[39966];
                
                r_data[39968] <= r_data[39967];
                
                r_data[39969] <= r_data[39968];
                
                r_data[39970] <= r_data[39969];
                
                r_data[39971] <= r_data[39970];
                
                r_data[39972] <= r_data[39971];
                
                r_data[39973] <= r_data[39972];
                
                r_data[39974] <= r_data[39973];
                
                r_data[39975] <= r_data[39974];
                
                r_data[39976] <= r_data[39975];
                
                r_data[39977] <= r_data[39976];
                
                r_data[39978] <= r_data[39977];
                
                r_data[39979] <= r_data[39978];
                
                r_data[39980] <= r_data[39979];
                
                r_data[39981] <= r_data[39980];
                
                r_data[39982] <= r_data[39981];
                
                r_data[39983] <= r_data[39982];
                
                r_data[39984] <= r_data[39983];
                
                r_data[39985] <= r_data[39984];
                
                r_data[39986] <= r_data[39985];
                
                r_data[39987] <= r_data[39986];
                
                r_data[39988] <= r_data[39987];
                
                r_data[39989] <= r_data[39988];
                
                r_data[39990] <= r_data[39989];
                
                r_data[39991] <= r_data[39990];
                
                r_data[39992] <= r_data[39991];
                
                r_data[39993] <= r_data[39992];
                
                r_data[39994] <= r_data[39993];
                
                r_data[39995] <= r_data[39994];
                
                r_data[39996] <= r_data[39995];
                
                r_data[39997] <= r_data[39996];
                
                r_data[39998] <= r_data[39997];
                
                r_data[39999] <= r_data[39998];
                
                r_data[40000] <= r_data[39999];
                
                r_data[40001] <= r_data[40000];
                
                r_data[40002] <= r_data[40001];
                
                r_data[40003] <= r_data[40002];
                
                r_data[40004] <= r_data[40003];
                
                r_data[40005] <= r_data[40004];
                
                r_data[40006] <= r_data[40005];
                
                r_data[40007] <= r_data[40006];
                
                r_data[40008] <= r_data[40007];
                
                r_data[40009] <= r_data[40008];
                
                r_data[40010] <= r_data[40009];
                
                r_data[40011] <= r_data[40010];
                
                r_data[40012] <= r_data[40011];
                
                r_data[40013] <= r_data[40012];
                
                r_data[40014] <= r_data[40013];
                
                r_data[40015] <= r_data[40014];
                
                r_data[40016] <= r_data[40015];
                
                r_data[40017] <= r_data[40016];
                
                r_data[40018] <= r_data[40017];
                
                r_data[40019] <= r_data[40018];
                
                r_data[40020] <= r_data[40019];
                
                r_data[40021] <= r_data[40020];
                
                r_data[40022] <= r_data[40021];
                
                r_data[40023] <= r_data[40022];
                
                r_data[40024] <= r_data[40023];
                
                r_data[40025] <= r_data[40024];
                
                r_data[40026] <= r_data[40025];
                
                r_data[40027] <= r_data[40026];
                
                r_data[40028] <= r_data[40027];
                
                r_data[40029] <= r_data[40028];
                
                r_data[40030] <= r_data[40029];
                
                r_data[40031] <= r_data[40030];
                
                r_data[40032] <= r_data[40031];
                
                r_data[40033] <= r_data[40032];
                
                r_data[40034] <= r_data[40033];
                
                r_data[40035] <= r_data[40034];
                
                r_data[40036] <= r_data[40035];
                
                r_data[40037] <= r_data[40036];
                
                r_data[40038] <= r_data[40037];
                
                r_data[40039] <= r_data[40038];
                
                r_data[40040] <= r_data[40039];
                
                r_data[40041] <= r_data[40040];
                
                r_data[40042] <= r_data[40041];
                
                r_data[40043] <= r_data[40042];
                
                r_data[40044] <= r_data[40043];
                
                r_data[40045] <= r_data[40044];
                
                r_data[40046] <= r_data[40045];
                
                r_data[40047] <= r_data[40046];
                
                r_data[40048] <= r_data[40047];
                
                r_data[40049] <= r_data[40048];
                
                r_data[40050] <= r_data[40049];
                
                r_data[40051] <= r_data[40050];
                
                r_data[40052] <= r_data[40051];
                
                r_data[40053] <= r_data[40052];
                
                r_data[40054] <= r_data[40053];
                
                r_data[40055] <= r_data[40054];
                
                r_data[40056] <= r_data[40055];
                
                r_data[40057] <= r_data[40056];
                
                r_data[40058] <= r_data[40057];
                
                r_data[40059] <= r_data[40058];
                
                r_data[40060] <= r_data[40059];
                
                r_data[40061] <= r_data[40060];
                
                r_data[40062] <= r_data[40061];
                
                r_data[40063] <= r_data[40062];
                
                r_data[40064] <= r_data[40063];
                
                r_data[40065] <= r_data[40064];
                
                r_data[40066] <= r_data[40065];
                
                r_data[40067] <= r_data[40066];
                
                r_data[40068] <= r_data[40067];
                
                r_data[40069] <= r_data[40068];
                
                r_data[40070] <= r_data[40069];
                
                r_data[40071] <= r_data[40070];
                
                r_data[40072] <= r_data[40071];
                
                r_data[40073] <= r_data[40072];
                
                r_data[40074] <= r_data[40073];
                
                r_data[40075] <= r_data[40074];
                
                r_data[40076] <= r_data[40075];
                
                r_data[40077] <= r_data[40076];
                
                r_data[40078] <= r_data[40077];
                
                r_data[40079] <= r_data[40078];
                
                r_data[40080] <= r_data[40079];
                
                r_data[40081] <= r_data[40080];
                
                r_data[40082] <= r_data[40081];
                
                r_data[40083] <= r_data[40082];
                
                r_data[40084] <= r_data[40083];
                
                r_data[40085] <= r_data[40084];
                
                r_data[40086] <= r_data[40085];
                
                r_data[40087] <= r_data[40086];
                
                r_data[40088] <= r_data[40087];
                
                r_data[40089] <= r_data[40088];
                
                r_data[40090] <= r_data[40089];
                
                r_data[40091] <= r_data[40090];
                
                r_data[40092] <= r_data[40091];
                
                r_data[40093] <= r_data[40092];
                
                r_data[40094] <= r_data[40093];
                
                r_data[40095] <= r_data[40094];
                
                r_data[40096] <= r_data[40095];
                
                r_data[40097] <= r_data[40096];
                
                r_data[40098] <= r_data[40097];
                
                r_data[40099] <= r_data[40098];
                
                r_data[40100] <= r_data[40099];
                
                r_data[40101] <= r_data[40100];
                
                r_data[40102] <= r_data[40101];
                
                r_data[40103] <= r_data[40102];
                
                r_data[40104] <= r_data[40103];
                
                r_data[40105] <= r_data[40104];
                
                r_data[40106] <= r_data[40105];
                
                r_data[40107] <= r_data[40106];
                
                r_data[40108] <= r_data[40107];
                
                r_data[40109] <= r_data[40108];
                
                r_data[40110] <= r_data[40109];
                
                r_data[40111] <= r_data[40110];
                
                r_data[40112] <= r_data[40111];
                
                r_data[40113] <= r_data[40112];
                
                r_data[40114] <= r_data[40113];
                
                r_data[40115] <= r_data[40114];
                
                r_data[40116] <= r_data[40115];
                
                r_data[40117] <= r_data[40116];
                
                r_data[40118] <= r_data[40117];
                
                r_data[40119] <= r_data[40118];
                
                r_data[40120] <= r_data[40119];
                
                r_data[40121] <= r_data[40120];
                
                r_data[40122] <= r_data[40121];
                
                r_data[40123] <= r_data[40122];
                
                r_data[40124] <= r_data[40123];
                
                r_data[40125] <= r_data[40124];
                
                r_data[40126] <= r_data[40125];
                
                r_data[40127] <= r_data[40126];
                
                r_data[40128] <= r_data[40127];
                
                r_data[40129] <= r_data[40128];
                
                r_data[40130] <= r_data[40129];
                
                r_data[40131] <= r_data[40130];
                
                r_data[40132] <= r_data[40131];
                
                r_data[40133] <= r_data[40132];
                
                r_data[40134] <= r_data[40133];
                
                r_data[40135] <= r_data[40134];
                
                r_data[40136] <= r_data[40135];
                
                r_data[40137] <= r_data[40136];
                
                r_data[40138] <= r_data[40137];
                
                r_data[40139] <= r_data[40138];
                
                r_data[40140] <= r_data[40139];
                
                r_data[40141] <= r_data[40140];
                
                r_data[40142] <= r_data[40141];
                
                r_data[40143] <= r_data[40142];
                
                r_data[40144] <= r_data[40143];
                
                r_data[40145] <= r_data[40144];
                
                r_data[40146] <= r_data[40145];
                
                r_data[40147] <= r_data[40146];
                
                r_data[40148] <= r_data[40147];
                
                r_data[40149] <= r_data[40148];
                
                r_data[40150] <= r_data[40149];
                
                r_data[40151] <= r_data[40150];
                
                r_data[40152] <= r_data[40151];
                
                r_data[40153] <= r_data[40152];
                
                r_data[40154] <= r_data[40153];
                
                r_data[40155] <= r_data[40154];
                
                r_data[40156] <= r_data[40155];
                
                r_data[40157] <= r_data[40156];
                
                r_data[40158] <= r_data[40157];
                
                r_data[40159] <= r_data[40158];
                
                r_data[40160] <= r_data[40159];
                
                r_data[40161] <= r_data[40160];
                
                r_data[40162] <= r_data[40161];
                
                r_data[40163] <= r_data[40162];
                
                r_data[40164] <= r_data[40163];
                
                r_data[40165] <= r_data[40164];
                
                r_data[40166] <= r_data[40165];
                
                r_data[40167] <= r_data[40166];
                
                r_data[40168] <= r_data[40167];
                
                r_data[40169] <= r_data[40168];
                
                r_data[40170] <= r_data[40169];
                
                r_data[40171] <= r_data[40170];
                
                r_data[40172] <= r_data[40171];
                
                r_data[40173] <= r_data[40172];
                
                r_data[40174] <= r_data[40173];
                
                r_data[40175] <= r_data[40174];
                
                r_data[40176] <= r_data[40175];
                
                r_data[40177] <= r_data[40176];
                
                r_data[40178] <= r_data[40177];
                
                r_data[40179] <= r_data[40178];
                
                r_data[40180] <= r_data[40179];
                
                r_data[40181] <= r_data[40180];
                
                r_data[40182] <= r_data[40181];
                
                r_data[40183] <= r_data[40182];
                
                r_data[40184] <= r_data[40183];
                
                r_data[40185] <= r_data[40184];
                
                r_data[40186] <= r_data[40185];
                
                r_data[40187] <= r_data[40186];
                
                r_data[40188] <= r_data[40187];
                
                r_data[40189] <= r_data[40188];
                
                r_data[40190] <= r_data[40189];
                
                r_data[40191] <= r_data[40190];
                
                r_data[40192] <= r_data[40191];
                
                r_data[40193] <= r_data[40192];
                
                r_data[40194] <= r_data[40193];
                
                r_data[40195] <= r_data[40194];
                
                r_data[40196] <= r_data[40195];
                
                r_data[40197] <= r_data[40196];
                
                r_data[40198] <= r_data[40197];
                
                r_data[40199] <= r_data[40198];
                
                r_data[40200] <= r_data[40199];
                
                r_data[40201] <= r_data[40200];
                
                r_data[40202] <= r_data[40201];
                
                r_data[40203] <= r_data[40202];
                
                r_data[40204] <= r_data[40203];
                
                r_data[40205] <= r_data[40204];
                
                r_data[40206] <= r_data[40205];
                
                r_data[40207] <= r_data[40206];
                
                r_data[40208] <= r_data[40207];
                
                r_data[40209] <= r_data[40208];
                
                r_data[40210] <= r_data[40209];
                
                r_data[40211] <= r_data[40210];
                
                r_data[40212] <= r_data[40211];
                
                r_data[40213] <= r_data[40212];
                
                r_data[40214] <= r_data[40213];
                
                r_data[40215] <= r_data[40214];
                
                r_data[40216] <= r_data[40215];
                
                r_data[40217] <= r_data[40216];
                
                r_data[40218] <= r_data[40217];
                
                r_data[40219] <= r_data[40218];
                
                r_data[40220] <= r_data[40219];
                
                r_data[40221] <= r_data[40220];
                
                r_data[40222] <= r_data[40221];
                
                r_data[40223] <= r_data[40222];
                
                r_data[40224] <= r_data[40223];
                
                r_data[40225] <= r_data[40224];
                
                r_data[40226] <= r_data[40225];
                
                r_data[40227] <= r_data[40226];
                
                r_data[40228] <= r_data[40227];
                
                r_data[40229] <= r_data[40228];
                
                r_data[40230] <= r_data[40229];
                
                r_data[40231] <= r_data[40230];
                
                r_data[40232] <= r_data[40231];
                
                r_data[40233] <= r_data[40232];
                
                r_data[40234] <= r_data[40233];
                
                r_data[40235] <= r_data[40234];
                
                r_data[40236] <= r_data[40235];
                
                r_data[40237] <= r_data[40236];
                
                r_data[40238] <= r_data[40237];
                
                r_data[40239] <= r_data[40238];
                
                r_data[40240] <= r_data[40239];
                
                r_data[40241] <= r_data[40240];
                
                r_data[40242] <= r_data[40241];
                
                r_data[40243] <= r_data[40242];
                
                r_data[40244] <= r_data[40243];
                
                r_data[40245] <= r_data[40244];
                
                r_data[40246] <= r_data[40245];
                
                r_data[40247] <= r_data[40246];
                
                r_data[40248] <= r_data[40247];
                
                r_data[40249] <= r_data[40248];
                
                r_data[40250] <= r_data[40249];
                
                r_data[40251] <= r_data[40250];
                
                r_data[40252] <= r_data[40251];
                
                r_data[40253] <= r_data[40252];
                
                r_data[40254] <= r_data[40253];
                
                r_data[40255] <= r_data[40254];
                
                r_data[40256] <= r_data[40255];
                
                r_data[40257] <= r_data[40256];
                
                r_data[40258] <= r_data[40257];
                
                r_data[40259] <= r_data[40258];
                
                r_data[40260] <= r_data[40259];
                
                r_data[40261] <= r_data[40260];
                
                r_data[40262] <= r_data[40261];
                
                r_data[40263] <= r_data[40262];
                
                r_data[40264] <= r_data[40263];
                
                r_data[40265] <= r_data[40264];
                
                r_data[40266] <= r_data[40265];
                
                r_data[40267] <= r_data[40266];
                
                r_data[40268] <= r_data[40267];
                
                r_data[40269] <= r_data[40268];
                
                r_data[40270] <= r_data[40269];
                
                r_data[40271] <= r_data[40270];
                
                r_data[40272] <= r_data[40271];
                
                r_data[40273] <= r_data[40272];
                
                r_data[40274] <= r_data[40273];
                
                r_data[40275] <= r_data[40274];
                
                r_data[40276] <= r_data[40275];
                
                r_data[40277] <= r_data[40276];
                
                r_data[40278] <= r_data[40277];
                
                r_data[40279] <= r_data[40278];
                
                r_data[40280] <= r_data[40279];
                
                r_data[40281] <= r_data[40280];
                
                r_data[40282] <= r_data[40281];
                
                r_data[40283] <= r_data[40282];
                
                r_data[40284] <= r_data[40283];
                
                r_data[40285] <= r_data[40284];
                
                r_data[40286] <= r_data[40285];
                
                r_data[40287] <= r_data[40286];
                
                r_data[40288] <= r_data[40287];
                
                r_data[40289] <= r_data[40288];
                
                r_data[40290] <= r_data[40289];
                
                r_data[40291] <= r_data[40290];
                
                r_data[40292] <= r_data[40291];
                
                r_data[40293] <= r_data[40292];
                
                r_data[40294] <= r_data[40293];
                
                r_data[40295] <= r_data[40294];
                
                r_data[40296] <= r_data[40295];
                
                r_data[40297] <= r_data[40296];
                
                r_data[40298] <= r_data[40297];
                
                r_data[40299] <= r_data[40298];
                
                r_data[40300] <= r_data[40299];
                
                r_data[40301] <= r_data[40300];
                
                r_data[40302] <= r_data[40301];
                
                r_data[40303] <= r_data[40302];
                
                r_data[40304] <= r_data[40303];
                
                r_data[40305] <= r_data[40304];
                
                r_data[40306] <= r_data[40305];
                
                r_data[40307] <= r_data[40306];
                
                r_data[40308] <= r_data[40307];
                
                r_data[40309] <= r_data[40308];
                
                r_data[40310] <= r_data[40309];
                
                r_data[40311] <= r_data[40310];
                
                r_data[40312] <= r_data[40311];
                
                r_data[40313] <= r_data[40312];
                
                r_data[40314] <= r_data[40313];
                
                r_data[40315] <= r_data[40314];
                
                r_data[40316] <= r_data[40315];
                
                r_data[40317] <= r_data[40316];
                
                r_data[40318] <= r_data[40317];
                
                r_data[40319] <= r_data[40318];
                
                r_data[40320] <= r_data[40319];
                
                r_data[40321] <= r_data[40320];
                
                r_data[40322] <= r_data[40321];
                
                r_data[40323] <= r_data[40322];
                
                r_data[40324] <= r_data[40323];
                
                r_data[40325] <= r_data[40324];
                
                r_data[40326] <= r_data[40325];
                
                r_data[40327] <= r_data[40326];
                
                r_data[40328] <= r_data[40327];
                
                r_data[40329] <= r_data[40328];
                
                r_data[40330] <= r_data[40329];
                
                r_data[40331] <= r_data[40330];
                
                r_data[40332] <= r_data[40331];
                
                r_data[40333] <= r_data[40332];
                
                r_data[40334] <= r_data[40333];
                
                r_data[40335] <= r_data[40334];
                
                r_data[40336] <= r_data[40335];
                
                r_data[40337] <= r_data[40336];
                
                r_data[40338] <= r_data[40337];
                
                r_data[40339] <= r_data[40338];
                
                r_data[40340] <= r_data[40339];
                
                r_data[40341] <= r_data[40340];
                
                r_data[40342] <= r_data[40341];
                
                r_data[40343] <= r_data[40342];
                
                r_data[40344] <= r_data[40343];
                
                r_data[40345] <= r_data[40344];
                
                r_data[40346] <= r_data[40345];
                
                r_data[40347] <= r_data[40346];
                
                r_data[40348] <= r_data[40347];
                
                r_data[40349] <= r_data[40348];
                
                r_data[40350] <= r_data[40349];
                
                r_data[40351] <= r_data[40350];
                
                r_data[40352] <= r_data[40351];
                
                r_data[40353] <= r_data[40352];
                
                r_data[40354] <= r_data[40353];
                
                r_data[40355] <= r_data[40354];
                
                r_data[40356] <= r_data[40355];
                
                r_data[40357] <= r_data[40356];
                
                r_data[40358] <= r_data[40357];
                
                r_data[40359] <= r_data[40358];
                
                r_data[40360] <= r_data[40359];
                
                r_data[40361] <= r_data[40360];
                
                r_data[40362] <= r_data[40361];
                
                r_data[40363] <= r_data[40362];
                
                r_data[40364] <= r_data[40363];
                
                r_data[40365] <= r_data[40364];
                
                r_data[40366] <= r_data[40365];
                
                r_data[40367] <= r_data[40366];
                
                r_data[40368] <= r_data[40367];
                
                r_data[40369] <= r_data[40368];
                
                r_data[40370] <= r_data[40369];
                
                r_data[40371] <= r_data[40370];
                
                r_data[40372] <= r_data[40371];
                
                r_data[40373] <= r_data[40372];
                
                r_data[40374] <= r_data[40373];
                
                r_data[40375] <= r_data[40374];
                
                r_data[40376] <= r_data[40375];
                
                r_data[40377] <= r_data[40376];
                
                r_data[40378] <= r_data[40377];
                
                r_data[40379] <= r_data[40378];
                
                r_data[40380] <= r_data[40379];
                
                r_data[40381] <= r_data[40380];
                
                r_data[40382] <= r_data[40381];
                
                r_data[40383] <= r_data[40382];
                
                r_data[40384] <= r_data[40383];
                
                r_data[40385] <= r_data[40384];
                
                r_data[40386] <= r_data[40385];
                
                r_data[40387] <= r_data[40386];
                
                r_data[40388] <= r_data[40387];
                
                r_data[40389] <= r_data[40388];
                
                r_data[40390] <= r_data[40389];
                
                r_data[40391] <= r_data[40390];
                
                r_data[40392] <= r_data[40391];
                
                r_data[40393] <= r_data[40392];
                
                r_data[40394] <= r_data[40393];
                
                r_data[40395] <= r_data[40394];
                
                r_data[40396] <= r_data[40395];
                
                r_data[40397] <= r_data[40396];
                
                r_data[40398] <= r_data[40397];
                
                r_data[40399] <= r_data[40398];
                
                r_data[40400] <= r_data[40399];
                
                r_data[40401] <= r_data[40400];
                
                r_data[40402] <= r_data[40401];
                
                r_data[40403] <= r_data[40402];
                
                r_data[40404] <= r_data[40403];
                
                r_data[40405] <= r_data[40404];
                
                r_data[40406] <= r_data[40405];
                
                r_data[40407] <= r_data[40406];
                
                r_data[40408] <= r_data[40407];
                
                r_data[40409] <= r_data[40408];
                
                r_data[40410] <= r_data[40409];
                
                r_data[40411] <= r_data[40410];
                
                r_data[40412] <= r_data[40411];
                
                r_data[40413] <= r_data[40412];
                
                r_data[40414] <= r_data[40413];
                
                r_data[40415] <= r_data[40414];
                
                r_data[40416] <= r_data[40415];
                
                r_data[40417] <= r_data[40416];
                
                r_data[40418] <= r_data[40417];
                
                r_data[40419] <= r_data[40418];
                
                r_data[40420] <= r_data[40419];
                
                r_data[40421] <= r_data[40420];
                
                r_data[40422] <= r_data[40421];
                
                r_data[40423] <= r_data[40422];
                
                r_data[40424] <= r_data[40423];
                
                r_data[40425] <= r_data[40424];
                
                r_data[40426] <= r_data[40425];
                
                r_data[40427] <= r_data[40426];
                
                r_data[40428] <= r_data[40427];
                
                r_data[40429] <= r_data[40428];
                
                r_data[40430] <= r_data[40429];
                
                r_data[40431] <= r_data[40430];
                
                r_data[40432] <= r_data[40431];
                
                r_data[40433] <= r_data[40432];
                
                r_data[40434] <= r_data[40433];
                
                r_data[40435] <= r_data[40434];
                
                r_data[40436] <= r_data[40435];
                
                r_data[40437] <= r_data[40436];
                
                r_data[40438] <= r_data[40437];
                
                r_data[40439] <= r_data[40438];
                
                r_data[40440] <= r_data[40439];
                
                r_data[40441] <= r_data[40440];
                
                r_data[40442] <= r_data[40441];
                
                r_data[40443] <= r_data[40442];
                
                r_data[40444] <= r_data[40443];
                
                r_data[40445] <= r_data[40444];
                
                r_data[40446] <= r_data[40445];
                
                r_data[40447] <= r_data[40446];
                
                r_data[40448] <= r_data[40447];
                
                r_data[40449] <= r_data[40448];
                
                r_data[40450] <= r_data[40449];
                
                r_data[40451] <= r_data[40450];
                
                r_data[40452] <= r_data[40451];
                
                r_data[40453] <= r_data[40452];
                
                r_data[40454] <= r_data[40453];
                
                r_data[40455] <= r_data[40454];
                
                r_data[40456] <= r_data[40455];
                
                r_data[40457] <= r_data[40456];
                
                r_data[40458] <= r_data[40457];
                
                r_data[40459] <= r_data[40458];
                
                r_data[40460] <= r_data[40459];
                
                r_data[40461] <= r_data[40460];
                
                r_data[40462] <= r_data[40461];
                
                r_data[40463] <= r_data[40462];
                
                r_data[40464] <= r_data[40463];
                
                r_data[40465] <= r_data[40464];
                
                r_data[40466] <= r_data[40465];
                
                r_data[40467] <= r_data[40466];
                
                r_data[40468] <= r_data[40467];
                
                r_data[40469] <= r_data[40468];
                
                r_data[40470] <= r_data[40469];
                
                r_data[40471] <= r_data[40470];
                
                r_data[40472] <= r_data[40471];
                
                r_data[40473] <= r_data[40472];
                
                r_data[40474] <= r_data[40473];
                
                r_data[40475] <= r_data[40474];
                
                r_data[40476] <= r_data[40475];
                
                r_data[40477] <= r_data[40476];
                
                r_data[40478] <= r_data[40477];
                
                r_data[40479] <= r_data[40478];
                
                r_data[40480] <= r_data[40479];
                
                r_data[40481] <= r_data[40480];
                
                r_data[40482] <= r_data[40481];
                
                r_data[40483] <= r_data[40482];
                
                r_data[40484] <= r_data[40483];
                
                r_data[40485] <= r_data[40484];
                
                r_data[40486] <= r_data[40485];
                
                r_data[40487] <= r_data[40486];
                
                r_data[40488] <= r_data[40487];
                
                r_data[40489] <= r_data[40488];
                
                r_data[40490] <= r_data[40489];
                
                r_data[40491] <= r_data[40490];
                
                r_data[40492] <= r_data[40491];
                
                r_data[40493] <= r_data[40492];
                
                r_data[40494] <= r_data[40493];
                
                r_data[40495] <= r_data[40494];
                
                r_data[40496] <= r_data[40495];
                
                r_data[40497] <= r_data[40496];
                
                r_data[40498] <= r_data[40497];
                
                r_data[40499] <= r_data[40498];
                
                r_data[40500] <= r_data[40499];
                
                r_data[40501] <= r_data[40500];
                
                r_data[40502] <= r_data[40501];
                
                r_data[40503] <= r_data[40502];
                
                r_data[40504] <= r_data[40503];
                
                r_data[40505] <= r_data[40504];
                
                r_data[40506] <= r_data[40505];
                
                r_data[40507] <= r_data[40506];
                
                r_data[40508] <= r_data[40507];
                
                r_data[40509] <= r_data[40508];
                
                r_data[40510] <= r_data[40509];
                
                r_data[40511] <= r_data[40510];
                
                r_data[40512] <= r_data[40511];
                
                r_data[40513] <= r_data[40512];
                
                r_data[40514] <= r_data[40513];
                
                r_data[40515] <= r_data[40514];
                
                r_data[40516] <= r_data[40515];
                
                r_data[40517] <= r_data[40516];
                
                r_data[40518] <= r_data[40517];
                
                r_data[40519] <= r_data[40518];
                
                r_data[40520] <= r_data[40519];
                
                r_data[40521] <= r_data[40520];
                
                r_data[40522] <= r_data[40521];
                
                r_data[40523] <= r_data[40522];
                
                r_data[40524] <= r_data[40523];
                
                r_data[40525] <= r_data[40524];
                
                r_data[40526] <= r_data[40525];
                
                r_data[40527] <= r_data[40526];
                
                r_data[40528] <= r_data[40527];
                
                r_data[40529] <= r_data[40528];
                
                r_data[40530] <= r_data[40529];
                
                r_data[40531] <= r_data[40530];
                
                r_data[40532] <= r_data[40531];
                
                r_data[40533] <= r_data[40532];
                
                r_data[40534] <= r_data[40533];
                
                r_data[40535] <= r_data[40534];
                
                r_data[40536] <= r_data[40535];
                
                r_data[40537] <= r_data[40536];
                
                r_data[40538] <= r_data[40537];
                
                r_data[40539] <= r_data[40538];
                
                r_data[40540] <= r_data[40539];
                
                r_data[40541] <= r_data[40540];
                
                r_data[40542] <= r_data[40541];
                
                r_data[40543] <= r_data[40542];
                
                r_data[40544] <= r_data[40543];
                
                r_data[40545] <= r_data[40544];
                
                r_data[40546] <= r_data[40545];
                
                r_data[40547] <= r_data[40546];
                
                r_data[40548] <= r_data[40547];
                
                r_data[40549] <= r_data[40548];
                
                r_data[40550] <= r_data[40549];
                
                r_data[40551] <= r_data[40550];
                
                r_data[40552] <= r_data[40551];
                
                r_data[40553] <= r_data[40552];
                
                r_data[40554] <= r_data[40553];
                
                r_data[40555] <= r_data[40554];
                
                r_data[40556] <= r_data[40555];
                
                r_data[40557] <= r_data[40556];
                
                r_data[40558] <= r_data[40557];
                
                r_data[40559] <= r_data[40558];
                
                r_data[40560] <= r_data[40559];
                
                r_data[40561] <= r_data[40560];
                
                r_data[40562] <= r_data[40561];
                
                r_data[40563] <= r_data[40562];
                
                r_data[40564] <= r_data[40563];
                
                r_data[40565] <= r_data[40564];
                
                r_data[40566] <= r_data[40565];
                
                r_data[40567] <= r_data[40566];
                
                r_data[40568] <= r_data[40567];
                
                r_data[40569] <= r_data[40568];
                
                r_data[40570] <= r_data[40569];
                
                r_data[40571] <= r_data[40570];
                
                r_data[40572] <= r_data[40571];
                
                r_data[40573] <= r_data[40572];
                
                r_data[40574] <= r_data[40573];
                
                r_data[40575] <= r_data[40574];
                
                r_data[40576] <= r_data[40575];
                
                r_data[40577] <= r_data[40576];
                
                r_data[40578] <= r_data[40577];
                
                r_data[40579] <= r_data[40578];
                
                r_data[40580] <= r_data[40579];
                
                r_data[40581] <= r_data[40580];
                
                r_data[40582] <= r_data[40581];
                
                r_data[40583] <= r_data[40582];
                
                r_data[40584] <= r_data[40583];
                
                r_data[40585] <= r_data[40584];
                
                r_data[40586] <= r_data[40585];
                
                r_data[40587] <= r_data[40586];
                
                r_data[40588] <= r_data[40587];
                
                r_data[40589] <= r_data[40588];
                
                r_data[40590] <= r_data[40589];
                
                r_data[40591] <= r_data[40590];
                
                r_data[40592] <= r_data[40591];
                
                r_data[40593] <= r_data[40592];
                
                r_data[40594] <= r_data[40593];
                
                r_data[40595] <= r_data[40594];
                
                r_data[40596] <= r_data[40595];
                
                r_data[40597] <= r_data[40596];
                
                r_data[40598] <= r_data[40597];
                
                r_data[40599] <= r_data[40598];
                
                r_data[40600] <= r_data[40599];
                
                r_data[40601] <= r_data[40600];
                
                r_data[40602] <= r_data[40601];
                
                r_data[40603] <= r_data[40602];
                
                r_data[40604] <= r_data[40603];
                
                r_data[40605] <= r_data[40604];
                
                r_data[40606] <= r_data[40605];
                
                r_data[40607] <= r_data[40606];
                
                r_data[40608] <= r_data[40607];
                
                r_data[40609] <= r_data[40608];
                
                r_data[40610] <= r_data[40609];
                
                r_data[40611] <= r_data[40610];
                
                r_data[40612] <= r_data[40611];
                
                r_data[40613] <= r_data[40612];
                
                r_data[40614] <= r_data[40613];
                
                r_data[40615] <= r_data[40614];
                
                r_data[40616] <= r_data[40615];
                
                r_data[40617] <= r_data[40616];
                
                r_data[40618] <= r_data[40617];
                
                r_data[40619] <= r_data[40618];
                
                r_data[40620] <= r_data[40619];
                
                r_data[40621] <= r_data[40620];
                
                r_data[40622] <= r_data[40621];
                
                r_data[40623] <= r_data[40622];
                
                r_data[40624] <= r_data[40623];
                
                r_data[40625] <= r_data[40624];
                
                r_data[40626] <= r_data[40625];
                
                r_data[40627] <= r_data[40626];
                
                r_data[40628] <= r_data[40627];
                
                r_data[40629] <= r_data[40628];
                
                r_data[40630] <= r_data[40629];
                
                r_data[40631] <= r_data[40630];
                
                r_data[40632] <= r_data[40631];
                
                r_data[40633] <= r_data[40632];
                
                r_data[40634] <= r_data[40633];
                
                r_data[40635] <= r_data[40634];
                
                r_data[40636] <= r_data[40635];
                
                r_data[40637] <= r_data[40636];
                
                r_data[40638] <= r_data[40637];
                
                r_data[40639] <= r_data[40638];
                
                r_data[40640] <= r_data[40639];
                
                r_data[40641] <= r_data[40640];
                
                r_data[40642] <= r_data[40641];
                
                r_data[40643] <= r_data[40642];
                
                r_data[40644] <= r_data[40643];
                
                r_data[40645] <= r_data[40644];
                
                r_data[40646] <= r_data[40645];
                
                r_data[40647] <= r_data[40646];
                
                r_data[40648] <= r_data[40647];
                
                r_data[40649] <= r_data[40648];
                
                r_data[40650] <= r_data[40649];
                
                r_data[40651] <= r_data[40650];
                
                r_data[40652] <= r_data[40651];
                
                r_data[40653] <= r_data[40652];
                
                r_data[40654] <= r_data[40653];
                
                r_data[40655] <= r_data[40654];
                
                r_data[40656] <= r_data[40655];
                
                r_data[40657] <= r_data[40656];
                
                r_data[40658] <= r_data[40657];
                
                r_data[40659] <= r_data[40658];
                
                r_data[40660] <= r_data[40659];
                
                r_data[40661] <= r_data[40660];
                
                r_data[40662] <= r_data[40661];
                
                r_data[40663] <= r_data[40662];
                
                r_data[40664] <= r_data[40663];
                
                r_data[40665] <= r_data[40664];
                
                r_data[40666] <= r_data[40665];
                
                r_data[40667] <= r_data[40666];
                
                r_data[40668] <= r_data[40667];
                
                r_data[40669] <= r_data[40668];
                
                r_data[40670] <= r_data[40669];
                
                r_data[40671] <= r_data[40670];
                
                r_data[40672] <= r_data[40671];
                
                r_data[40673] <= r_data[40672];
                
                r_data[40674] <= r_data[40673];
                
                r_data[40675] <= r_data[40674];
                
                r_data[40676] <= r_data[40675];
                
                r_data[40677] <= r_data[40676];
                
                r_data[40678] <= r_data[40677];
                
                r_data[40679] <= r_data[40678];
                
                r_data[40680] <= r_data[40679];
                
                r_data[40681] <= r_data[40680];
                
                r_data[40682] <= r_data[40681];
                
                r_data[40683] <= r_data[40682];
                
                r_data[40684] <= r_data[40683];
                
                r_data[40685] <= r_data[40684];
                
                r_data[40686] <= r_data[40685];
                
                r_data[40687] <= r_data[40686];
                
                r_data[40688] <= r_data[40687];
                
                r_data[40689] <= r_data[40688];
                
                r_data[40690] <= r_data[40689];
                
                r_data[40691] <= r_data[40690];
                
                r_data[40692] <= r_data[40691];
                
                r_data[40693] <= r_data[40692];
                
                r_data[40694] <= r_data[40693];
                
                r_data[40695] <= r_data[40694];
                
                r_data[40696] <= r_data[40695];
                
                r_data[40697] <= r_data[40696];
                
                r_data[40698] <= r_data[40697];
                
                r_data[40699] <= r_data[40698];
                
                r_data[40700] <= r_data[40699];
                
                r_data[40701] <= r_data[40700];
                
                r_data[40702] <= r_data[40701];
                
                r_data[40703] <= r_data[40702];
                
                r_data[40704] <= r_data[40703];
                
                r_data[40705] <= r_data[40704];
                
                r_data[40706] <= r_data[40705];
                
                r_data[40707] <= r_data[40706];
                
                r_data[40708] <= r_data[40707];
                
                r_data[40709] <= r_data[40708];
                
                r_data[40710] <= r_data[40709];
                
                r_data[40711] <= r_data[40710];
                
                r_data[40712] <= r_data[40711];
                
                r_data[40713] <= r_data[40712];
                
                r_data[40714] <= r_data[40713];
                
                r_data[40715] <= r_data[40714];
                
                r_data[40716] <= r_data[40715];
                
                r_data[40717] <= r_data[40716];
                
                r_data[40718] <= r_data[40717];
                
                r_data[40719] <= r_data[40718];
                
                r_data[40720] <= r_data[40719];
                
                r_data[40721] <= r_data[40720];
                
                r_data[40722] <= r_data[40721];
                
                r_data[40723] <= r_data[40722];
                
                r_data[40724] <= r_data[40723];
                
                r_data[40725] <= r_data[40724];
                
                r_data[40726] <= r_data[40725];
                
                r_data[40727] <= r_data[40726];
                
                r_data[40728] <= r_data[40727];
                
                r_data[40729] <= r_data[40728];
                
                r_data[40730] <= r_data[40729];
                
                r_data[40731] <= r_data[40730];
                
                r_data[40732] <= r_data[40731];
                
                r_data[40733] <= r_data[40732];
                
                r_data[40734] <= r_data[40733];
                
                r_data[40735] <= r_data[40734];
                
                r_data[40736] <= r_data[40735];
                
                r_data[40737] <= r_data[40736];
                
                r_data[40738] <= r_data[40737];
                
                r_data[40739] <= r_data[40738];
                
                r_data[40740] <= r_data[40739];
                
                r_data[40741] <= r_data[40740];
                
                r_data[40742] <= r_data[40741];
                
                r_data[40743] <= r_data[40742];
                
                r_data[40744] <= r_data[40743];
                
                r_data[40745] <= r_data[40744];
                
                r_data[40746] <= r_data[40745];
                
                r_data[40747] <= r_data[40746];
                
                r_data[40748] <= r_data[40747];
                
                r_data[40749] <= r_data[40748];
                
                r_data[40750] <= r_data[40749];
                
                r_data[40751] <= r_data[40750];
                
                r_data[40752] <= r_data[40751];
                
                r_data[40753] <= r_data[40752];
                
                r_data[40754] <= r_data[40753];
                
                r_data[40755] <= r_data[40754];
                
                r_data[40756] <= r_data[40755];
                
                r_data[40757] <= r_data[40756];
                
                r_data[40758] <= r_data[40757];
                
                r_data[40759] <= r_data[40758];
                
                r_data[40760] <= r_data[40759];
                
                r_data[40761] <= r_data[40760];
                
                r_data[40762] <= r_data[40761];
                
                r_data[40763] <= r_data[40762];
                
                r_data[40764] <= r_data[40763];
                
                r_data[40765] <= r_data[40764];
                
                r_data[40766] <= r_data[40765];
                
                r_data[40767] <= r_data[40766];
                
                r_data[40768] <= r_data[40767];
                
                r_data[40769] <= r_data[40768];
                
                r_data[40770] <= r_data[40769];
                
                r_data[40771] <= r_data[40770];
                
                r_data[40772] <= r_data[40771];
                
                r_data[40773] <= r_data[40772];
                
                r_data[40774] <= r_data[40773];
                
                r_data[40775] <= r_data[40774];
                
                r_data[40776] <= r_data[40775];
                
                r_data[40777] <= r_data[40776];
                
                r_data[40778] <= r_data[40777];
                
                r_data[40779] <= r_data[40778];
                
                r_data[40780] <= r_data[40779];
                
                r_data[40781] <= r_data[40780];
                
                r_data[40782] <= r_data[40781];
                
                r_data[40783] <= r_data[40782];
                
                r_data[40784] <= r_data[40783];
                
                r_data[40785] <= r_data[40784];
                
                r_data[40786] <= r_data[40785];
                
                r_data[40787] <= r_data[40786];
                
                r_data[40788] <= r_data[40787];
                
                r_data[40789] <= r_data[40788];
                
                r_data[40790] <= r_data[40789];
                
                r_data[40791] <= r_data[40790];
                
                r_data[40792] <= r_data[40791];
                
                r_data[40793] <= r_data[40792];
                
                r_data[40794] <= r_data[40793];
                
                r_data[40795] <= r_data[40794];
                
                r_data[40796] <= r_data[40795];
                
                r_data[40797] <= r_data[40796];
                
                r_data[40798] <= r_data[40797];
                
                r_data[40799] <= r_data[40798];
                
                r_data[40800] <= r_data[40799];
                
                r_data[40801] <= r_data[40800];
                
                r_data[40802] <= r_data[40801];
                
                r_data[40803] <= r_data[40802];
                
                r_data[40804] <= r_data[40803];
                
                r_data[40805] <= r_data[40804];
                
                r_data[40806] <= r_data[40805];
                
                r_data[40807] <= r_data[40806];
                
                r_data[40808] <= r_data[40807];
                
                r_data[40809] <= r_data[40808];
                
                r_data[40810] <= r_data[40809];
                
                r_data[40811] <= r_data[40810];
                
                r_data[40812] <= r_data[40811];
                
                r_data[40813] <= r_data[40812];
                
                r_data[40814] <= r_data[40813];
                
                r_data[40815] <= r_data[40814];
                
                r_data[40816] <= r_data[40815];
                
                r_data[40817] <= r_data[40816];
                
                r_data[40818] <= r_data[40817];
                
                r_data[40819] <= r_data[40818];
                
                r_data[40820] <= r_data[40819];
                
                r_data[40821] <= r_data[40820];
                
                r_data[40822] <= r_data[40821];
                
                r_data[40823] <= r_data[40822];
                
                r_data[40824] <= r_data[40823];
                
                r_data[40825] <= r_data[40824];
                
                r_data[40826] <= r_data[40825];
                
                r_data[40827] <= r_data[40826];
                
                r_data[40828] <= r_data[40827];
                
                r_data[40829] <= r_data[40828];
                
                r_data[40830] <= r_data[40829];
                
                r_data[40831] <= r_data[40830];
                
                r_data[40832] <= r_data[40831];
                
                r_data[40833] <= r_data[40832];
                
                r_data[40834] <= r_data[40833];
                
                r_data[40835] <= r_data[40834];
                
                r_data[40836] <= r_data[40835];
                
                r_data[40837] <= r_data[40836];
                
                r_data[40838] <= r_data[40837];
                
                r_data[40839] <= r_data[40838];
                
                r_data[40840] <= r_data[40839];
                
                r_data[40841] <= r_data[40840];
                
                r_data[40842] <= r_data[40841];
                
                r_data[40843] <= r_data[40842];
                
                r_data[40844] <= r_data[40843];
                
                r_data[40845] <= r_data[40844];
                
                r_data[40846] <= r_data[40845];
                
                r_data[40847] <= r_data[40846];
                
                r_data[40848] <= r_data[40847];
                
                r_data[40849] <= r_data[40848];
                
                r_data[40850] <= r_data[40849];
                
                r_data[40851] <= r_data[40850];
                
                r_data[40852] <= r_data[40851];
                
                r_data[40853] <= r_data[40852];
                
                r_data[40854] <= r_data[40853];
                
                r_data[40855] <= r_data[40854];
                
                r_data[40856] <= r_data[40855];
                
                r_data[40857] <= r_data[40856];
                
                r_data[40858] <= r_data[40857];
                
                r_data[40859] <= r_data[40858];
                
                r_data[40860] <= r_data[40859];
                
                r_data[40861] <= r_data[40860];
                
                r_data[40862] <= r_data[40861];
                
                r_data[40863] <= r_data[40862];
                
                r_data[40864] <= r_data[40863];
                
                r_data[40865] <= r_data[40864];
                
                r_data[40866] <= r_data[40865];
                
                r_data[40867] <= r_data[40866];
                
                r_data[40868] <= r_data[40867];
                
                r_data[40869] <= r_data[40868];
                
                r_data[40870] <= r_data[40869];
                
                r_data[40871] <= r_data[40870];
                
                r_data[40872] <= r_data[40871];
                
                r_data[40873] <= r_data[40872];
                
                r_data[40874] <= r_data[40873];
                
                r_data[40875] <= r_data[40874];
                
                r_data[40876] <= r_data[40875];
                
                r_data[40877] <= r_data[40876];
                
                r_data[40878] <= r_data[40877];
                
                r_data[40879] <= r_data[40878];
                
                r_data[40880] <= r_data[40879];
                
                r_data[40881] <= r_data[40880];
                
                r_data[40882] <= r_data[40881];
                
                r_data[40883] <= r_data[40882];
                
                r_data[40884] <= r_data[40883];
                
                r_data[40885] <= r_data[40884];
                
                r_data[40886] <= r_data[40885];
                
                r_data[40887] <= r_data[40886];
                
                r_data[40888] <= r_data[40887];
                
                r_data[40889] <= r_data[40888];
                
                r_data[40890] <= r_data[40889];
                
                r_data[40891] <= r_data[40890];
                
                r_data[40892] <= r_data[40891];
                
                r_data[40893] <= r_data[40892];
                
                r_data[40894] <= r_data[40893];
                
                r_data[40895] <= r_data[40894];
                
                r_data[40896] <= r_data[40895];
                
                r_data[40897] <= r_data[40896];
                
                r_data[40898] <= r_data[40897];
                
                r_data[40899] <= r_data[40898];
                
                r_data[40900] <= r_data[40899];
                
                r_data[40901] <= r_data[40900];
                
                r_data[40902] <= r_data[40901];
                
                r_data[40903] <= r_data[40902];
                
                r_data[40904] <= r_data[40903];
                
                r_data[40905] <= r_data[40904];
                
                r_data[40906] <= r_data[40905];
                
                r_data[40907] <= r_data[40906];
                
                r_data[40908] <= r_data[40907];
                
                r_data[40909] <= r_data[40908];
                
                r_data[40910] <= r_data[40909];
                
                r_data[40911] <= r_data[40910];
                
                r_data[40912] <= r_data[40911];
                
                r_data[40913] <= r_data[40912];
                
                r_data[40914] <= r_data[40913];
                
                r_data[40915] <= r_data[40914];
                
                r_data[40916] <= r_data[40915];
                
                r_data[40917] <= r_data[40916];
                
                r_data[40918] <= r_data[40917];
                
                r_data[40919] <= r_data[40918];
                
                r_data[40920] <= r_data[40919];
                
                r_data[40921] <= r_data[40920];
                
                r_data[40922] <= r_data[40921];
                
                r_data[40923] <= r_data[40922];
                
                r_data[40924] <= r_data[40923];
                
                r_data[40925] <= r_data[40924];
                
                r_data[40926] <= r_data[40925];
                
                r_data[40927] <= r_data[40926];
                
                r_data[40928] <= r_data[40927];
                
                r_data[40929] <= r_data[40928];
                
                r_data[40930] <= r_data[40929];
                
                r_data[40931] <= r_data[40930];
                
                r_data[40932] <= r_data[40931];
                
                r_data[40933] <= r_data[40932];
                
                r_data[40934] <= r_data[40933];
                
                r_data[40935] <= r_data[40934];
                
                r_data[40936] <= r_data[40935];
                
                r_data[40937] <= r_data[40936];
                
                r_data[40938] <= r_data[40937];
                
                r_data[40939] <= r_data[40938];
                
                r_data[40940] <= r_data[40939];
                
                r_data[40941] <= r_data[40940];
                
                r_data[40942] <= r_data[40941];
                
                r_data[40943] <= r_data[40942];
                
                r_data[40944] <= r_data[40943];
                
                r_data[40945] <= r_data[40944];
                
                r_data[40946] <= r_data[40945];
                
                r_data[40947] <= r_data[40946];
                
                r_data[40948] <= r_data[40947];
                
                r_data[40949] <= r_data[40948];
                
                r_data[40950] <= r_data[40949];
                
                r_data[40951] <= r_data[40950];
                
                r_data[40952] <= r_data[40951];
                
                r_data[40953] <= r_data[40952];
                
                r_data[40954] <= r_data[40953];
                
                r_data[40955] <= r_data[40954];
                
                r_data[40956] <= r_data[40955];
                
                r_data[40957] <= r_data[40956];
                
                r_data[40958] <= r_data[40957];
                
                r_data[40959] <= r_data[40958];
                
                r_data[40960] <= r_data[40959];
                
                r_data[40961] <= r_data[40960];
                
                r_data[40962] <= r_data[40961];
                
                r_data[40963] <= r_data[40962];
                
                r_data[40964] <= r_data[40963];
                
                r_data[40965] <= r_data[40964];
                
                r_data[40966] <= r_data[40965];
                
                r_data[40967] <= r_data[40966];
                
                r_data[40968] <= r_data[40967];
                
                r_data[40969] <= r_data[40968];
                
                r_data[40970] <= r_data[40969];
                
                r_data[40971] <= r_data[40970];
                
                r_data[40972] <= r_data[40971];
                
                r_data[40973] <= r_data[40972];
                
                r_data[40974] <= r_data[40973];
                
                r_data[40975] <= r_data[40974];
                
                r_data[40976] <= r_data[40975];
                
                r_data[40977] <= r_data[40976];
                
                r_data[40978] <= r_data[40977];
                
                r_data[40979] <= r_data[40978];
                
                r_data[40980] <= r_data[40979];
                
                r_data[40981] <= r_data[40980];
                
                r_data[40982] <= r_data[40981];
                
                r_data[40983] <= r_data[40982];
                
                r_data[40984] <= r_data[40983];
                
                r_data[40985] <= r_data[40984];
                
                r_data[40986] <= r_data[40985];
                
                r_data[40987] <= r_data[40986];
                
                r_data[40988] <= r_data[40987];
                
                r_data[40989] <= r_data[40988];
                
                r_data[40990] <= r_data[40989];
                
                r_data[40991] <= r_data[40990];
                
                r_data[40992] <= r_data[40991];
                
                r_data[40993] <= r_data[40992];
                
                r_data[40994] <= r_data[40993];
                
                r_data[40995] <= r_data[40994];
                
                r_data[40996] <= r_data[40995];
                
                r_data[40997] <= r_data[40996];
                
                r_data[40998] <= r_data[40997];
                
                r_data[40999] <= r_data[40998];
                
                r_data[41000] <= r_data[40999];
                
                r_data[41001] <= r_data[41000];
                
                r_data[41002] <= r_data[41001];
                
                r_data[41003] <= r_data[41002];
                
                r_data[41004] <= r_data[41003];
                
                r_data[41005] <= r_data[41004];
                
                r_data[41006] <= r_data[41005];
                
                r_data[41007] <= r_data[41006];
                
                r_data[41008] <= r_data[41007];
                
                r_data[41009] <= r_data[41008];
                
                r_data[41010] <= r_data[41009];
                
                r_data[41011] <= r_data[41010];
                
                r_data[41012] <= r_data[41011];
                
                r_data[41013] <= r_data[41012];
                
                r_data[41014] <= r_data[41013];
                
                r_data[41015] <= r_data[41014];
                
                r_data[41016] <= r_data[41015];
                
                r_data[41017] <= r_data[41016];
                
                r_data[41018] <= r_data[41017];
                
                r_data[41019] <= r_data[41018];
                
                r_data[41020] <= r_data[41019];
                
                r_data[41021] <= r_data[41020];
                
                r_data[41022] <= r_data[41021];
                
                r_data[41023] <= r_data[41022];
                
                r_data[41024] <= r_data[41023];
                
                r_data[41025] <= r_data[41024];
                
                r_data[41026] <= r_data[41025];
                
                r_data[41027] <= r_data[41026];
                
                r_data[41028] <= r_data[41027];
                
                r_data[41029] <= r_data[41028];
                
                r_data[41030] <= r_data[41029];
                
                r_data[41031] <= r_data[41030];
                
                r_data[41032] <= r_data[41031];
                
                r_data[41033] <= r_data[41032];
                
                r_data[41034] <= r_data[41033];
                
                r_data[41035] <= r_data[41034];
                
                r_data[41036] <= r_data[41035];
                
                r_data[41037] <= r_data[41036];
                
                r_data[41038] <= r_data[41037];
                
                r_data[41039] <= r_data[41038];
                
                r_data[41040] <= r_data[41039];
                
                r_data[41041] <= r_data[41040];
                
                r_data[41042] <= r_data[41041];
                
                r_data[41043] <= r_data[41042];
                
                r_data[41044] <= r_data[41043];
                
                r_data[41045] <= r_data[41044];
                
                r_data[41046] <= r_data[41045];
                
                r_data[41047] <= r_data[41046];
                
                r_data[41048] <= r_data[41047];
                
                r_data[41049] <= r_data[41048];
                
                r_data[41050] <= r_data[41049];
                
                r_data[41051] <= r_data[41050];
                
                r_data[41052] <= r_data[41051];
                
                r_data[41053] <= r_data[41052];
                
                r_data[41054] <= r_data[41053];
                
                r_data[41055] <= r_data[41054];
                
                r_data[41056] <= r_data[41055];
                
                r_data[41057] <= r_data[41056];
                
                r_data[41058] <= r_data[41057];
                
                r_data[41059] <= r_data[41058];
                
                r_data[41060] <= r_data[41059];
                
                r_data[41061] <= r_data[41060];
                
                r_data[41062] <= r_data[41061];
                
                r_data[41063] <= r_data[41062];
                
                r_data[41064] <= r_data[41063];
                
                r_data[41065] <= r_data[41064];
                
                r_data[41066] <= r_data[41065];
                
                r_data[41067] <= r_data[41066];
                
                r_data[41068] <= r_data[41067];
                
                r_data[41069] <= r_data[41068];
                
                r_data[41070] <= r_data[41069];
                
                r_data[41071] <= r_data[41070];
                
                r_data[41072] <= r_data[41071];
                
                r_data[41073] <= r_data[41072];
                
                r_data[41074] <= r_data[41073];
                
                r_data[41075] <= r_data[41074];
                
                r_data[41076] <= r_data[41075];
                
                r_data[41077] <= r_data[41076];
                
                r_data[41078] <= r_data[41077];
                
                r_data[41079] <= r_data[41078];
                
                r_data[41080] <= r_data[41079];
                
                r_data[41081] <= r_data[41080];
                
                r_data[41082] <= r_data[41081];
                
                r_data[41083] <= r_data[41082];
                
                r_data[41084] <= r_data[41083];
                
                r_data[41085] <= r_data[41084];
                
                r_data[41086] <= r_data[41085];
                
                r_data[41087] <= r_data[41086];
                
                r_data[41088] <= r_data[41087];
                
                r_data[41089] <= r_data[41088];
                
                r_data[41090] <= r_data[41089];
                
                r_data[41091] <= r_data[41090];
                
                r_data[41092] <= r_data[41091];
                
                r_data[41093] <= r_data[41092];
                
                r_data[41094] <= r_data[41093];
                
                r_data[41095] <= r_data[41094];
                
                r_data[41096] <= r_data[41095];
                
                r_data[41097] <= r_data[41096];
                
                r_data[41098] <= r_data[41097];
                
                r_data[41099] <= r_data[41098];
                
                r_data[41100] <= r_data[41099];
                
                r_data[41101] <= r_data[41100];
                
                r_data[41102] <= r_data[41101];
                
                r_data[41103] <= r_data[41102];
                
                r_data[41104] <= r_data[41103];
                
                r_data[41105] <= r_data[41104];
                
                r_data[41106] <= r_data[41105];
                
                r_data[41107] <= r_data[41106];
                
                r_data[41108] <= r_data[41107];
                
                r_data[41109] <= r_data[41108];
                
                r_data[41110] <= r_data[41109];
                
                r_data[41111] <= r_data[41110];
                
                r_data[41112] <= r_data[41111];
                
                r_data[41113] <= r_data[41112];
                
                r_data[41114] <= r_data[41113];
                
                r_data[41115] <= r_data[41114];
                
                r_data[41116] <= r_data[41115];
                
                r_data[41117] <= r_data[41116];
                
                r_data[41118] <= r_data[41117];
                
                r_data[41119] <= r_data[41118];
                
                r_data[41120] <= r_data[41119];
                
                r_data[41121] <= r_data[41120];
                
                r_data[41122] <= r_data[41121];
                
                r_data[41123] <= r_data[41122];
                
                r_data[41124] <= r_data[41123];
                
                r_data[41125] <= r_data[41124];
                
                r_data[41126] <= r_data[41125];
                
                r_data[41127] <= r_data[41126];
                
                r_data[41128] <= r_data[41127];
                
                r_data[41129] <= r_data[41128];
                
                r_data[41130] <= r_data[41129];
                
                r_data[41131] <= r_data[41130];
                
                r_data[41132] <= r_data[41131];
                
                r_data[41133] <= r_data[41132];
                
                r_data[41134] <= r_data[41133];
                
                r_data[41135] <= r_data[41134];
                
                r_data[41136] <= r_data[41135];
                
                r_data[41137] <= r_data[41136];
                
                r_data[41138] <= r_data[41137];
                
                r_data[41139] <= r_data[41138];
                
                r_data[41140] <= r_data[41139];
                
                r_data[41141] <= r_data[41140];
                
                r_data[41142] <= r_data[41141];
                
                r_data[41143] <= r_data[41142];
                
                r_data[41144] <= r_data[41143];
                
                r_data[41145] <= r_data[41144];
                
                r_data[41146] <= r_data[41145];
                
                r_data[41147] <= r_data[41146];
                
                r_data[41148] <= r_data[41147];
                
                r_data[41149] <= r_data[41148];
                
                r_data[41150] <= r_data[41149];
                
                r_data[41151] <= r_data[41150];
                
                r_data[41152] <= r_data[41151];
                
                r_data[41153] <= r_data[41152];
                
                r_data[41154] <= r_data[41153];
                
                r_data[41155] <= r_data[41154];
                
                r_data[41156] <= r_data[41155];
                
                r_data[41157] <= r_data[41156];
                
                r_data[41158] <= r_data[41157];
                
                r_data[41159] <= r_data[41158];
                
                r_data[41160] <= r_data[41159];
                
                r_data[41161] <= r_data[41160];
                
                r_data[41162] <= r_data[41161];
                
                r_data[41163] <= r_data[41162];
                
                r_data[41164] <= r_data[41163];
                
                r_data[41165] <= r_data[41164];
                
                r_data[41166] <= r_data[41165];
                
                r_data[41167] <= r_data[41166];
                
                r_data[41168] <= r_data[41167];
                
                r_data[41169] <= r_data[41168];
                
                r_data[41170] <= r_data[41169];
                
                r_data[41171] <= r_data[41170];
                
                r_data[41172] <= r_data[41171];
                
                r_data[41173] <= r_data[41172];
                
                r_data[41174] <= r_data[41173];
                
                r_data[41175] <= r_data[41174];
                
                r_data[41176] <= r_data[41175];
                
                r_data[41177] <= r_data[41176];
                
                r_data[41178] <= r_data[41177];
                
                r_data[41179] <= r_data[41178];
                
                r_data[41180] <= r_data[41179];
                
                r_data[41181] <= r_data[41180];
                
                r_data[41182] <= r_data[41181];
                
                r_data[41183] <= r_data[41182];
                
                r_data[41184] <= r_data[41183];
                
                r_data[41185] <= r_data[41184];
                
                r_data[41186] <= r_data[41185];
                
                r_data[41187] <= r_data[41186];
                
                r_data[41188] <= r_data[41187];
                
                r_data[41189] <= r_data[41188];
                
                r_data[41190] <= r_data[41189];
                
                r_data[41191] <= r_data[41190];
                
                r_data[41192] <= r_data[41191];
                
                r_data[41193] <= r_data[41192];
                
                r_data[41194] <= r_data[41193];
                
                r_data[41195] <= r_data[41194];
                
                r_data[41196] <= r_data[41195];
                
                r_data[41197] <= r_data[41196];
                
                r_data[41198] <= r_data[41197];
                
                r_data[41199] <= r_data[41198];
                
                r_data[41200] <= r_data[41199];
                
                r_data[41201] <= r_data[41200];
                
                r_data[41202] <= r_data[41201];
                
                r_data[41203] <= r_data[41202];
                
                r_data[41204] <= r_data[41203];
                
                r_data[41205] <= r_data[41204];
                
                r_data[41206] <= r_data[41205];
                
                r_data[41207] <= r_data[41206];
                
                r_data[41208] <= r_data[41207];
                
                r_data[41209] <= r_data[41208];
                
                r_data[41210] <= r_data[41209];
                
                r_data[41211] <= r_data[41210];
                
                r_data[41212] <= r_data[41211];
                
                r_data[41213] <= r_data[41212];
                
                r_data[41214] <= r_data[41213];
                
                r_data[41215] <= r_data[41214];
                
                r_data[41216] <= r_data[41215];
                
                r_data[41217] <= r_data[41216];
                
                r_data[41218] <= r_data[41217];
                
                r_data[41219] <= r_data[41218];
                
                r_data[41220] <= r_data[41219];
                
                r_data[41221] <= r_data[41220];
                
                r_data[41222] <= r_data[41221];
                
                r_data[41223] <= r_data[41222];
                
                r_data[41224] <= r_data[41223];
                
                r_data[41225] <= r_data[41224];
                
                r_data[41226] <= r_data[41225];
                
                r_data[41227] <= r_data[41226];
                
                r_data[41228] <= r_data[41227];
                
                r_data[41229] <= r_data[41228];
                
                r_data[41230] <= r_data[41229];
                
                r_data[41231] <= r_data[41230];
                
                r_data[41232] <= r_data[41231];
                
                r_data[41233] <= r_data[41232];
                
                r_data[41234] <= r_data[41233];
                
                r_data[41235] <= r_data[41234];
                
                r_data[41236] <= r_data[41235];
                
                r_data[41237] <= r_data[41236];
                
                r_data[41238] <= r_data[41237];
                
                r_data[41239] <= r_data[41238];
                
                r_data[41240] <= r_data[41239];
                
                r_data[41241] <= r_data[41240];
                
                r_data[41242] <= r_data[41241];
                
                r_data[41243] <= r_data[41242];
                
                r_data[41244] <= r_data[41243];
                
                r_data[41245] <= r_data[41244];
                
                r_data[41246] <= r_data[41245];
                
                r_data[41247] <= r_data[41246];
                
                r_data[41248] <= r_data[41247];
                
                r_data[41249] <= r_data[41248];
                
                r_data[41250] <= r_data[41249];
                
                r_data[41251] <= r_data[41250];
                
                r_data[41252] <= r_data[41251];
                
                r_data[41253] <= r_data[41252];
                
                r_data[41254] <= r_data[41253];
                
                r_data[41255] <= r_data[41254];
                
                r_data[41256] <= r_data[41255];
                
                r_data[41257] <= r_data[41256];
                
                r_data[41258] <= r_data[41257];
                
                r_data[41259] <= r_data[41258];
                
                r_data[41260] <= r_data[41259];
                
                r_data[41261] <= r_data[41260];
                
                r_data[41262] <= r_data[41261];
                
                r_data[41263] <= r_data[41262];
                
                r_data[41264] <= r_data[41263];
                
                r_data[41265] <= r_data[41264];
                
                r_data[41266] <= r_data[41265];
                
                r_data[41267] <= r_data[41266];
                
                r_data[41268] <= r_data[41267];
                
                r_data[41269] <= r_data[41268];
                
                r_data[41270] <= r_data[41269];
                
                r_data[41271] <= r_data[41270];
                
                r_data[41272] <= r_data[41271];
                
                r_data[41273] <= r_data[41272];
                
                r_data[41274] <= r_data[41273];
                
                r_data[41275] <= r_data[41274];
                
                r_data[41276] <= r_data[41275];
                
                r_data[41277] <= r_data[41276];
                
                r_data[41278] <= r_data[41277];
                
                r_data[41279] <= r_data[41278];
                
                r_data[41280] <= r_data[41279];
                
                r_data[41281] <= r_data[41280];
                
                r_data[41282] <= r_data[41281];
                
                r_data[41283] <= r_data[41282];
                
                r_data[41284] <= r_data[41283];
                
                r_data[41285] <= r_data[41284];
                
                r_data[41286] <= r_data[41285];
                
                r_data[41287] <= r_data[41286];
                
                r_data[41288] <= r_data[41287];
                
                r_data[41289] <= r_data[41288];
                
                r_data[41290] <= r_data[41289];
                
                r_data[41291] <= r_data[41290];
                
                r_data[41292] <= r_data[41291];
                
                r_data[41293] <= r_data[41292];
                
                r_data[41294] <= r_data[41293];
                
                r_data[41295] <= r_data[41294];
                
                r_data[41296] <= r_data[41295];
                
                r_data[41297] <= r_data[41296];
                
                r_data[41298] <= r_data[41297];
                
                r_data[41299] <= r_data[41298];
                
                r_data[41300] <= r_data[41299];
                
                r_data[41301] <= r_data[41300];
                
                r_data[41302] <= r_data[41301];
                
                r_data[41303] <= r_data[41302];
                
                r_data[41304] <= r_data[41303];
                
                r_data[41305] <= r_data[41304];
                
                r_data[41306] <= r_data[41305];
                
                r_data[41307] <= r_data[41306];
                
                r_data[41308] <= r_data[41307];
                
                r_data[41309] <= r_data[41308];
                
                r_data[41310] <= r_data[41309];
                
                r_data[41311] <= r_data[41310];
                
                r_data[41312] <= r_data[41311];
                
                r_data[41313] <= r_data[41312];
                
                r_data[41314] <= r_data[41313];
                
                r_data[41315] <= r_data[41314];
                
                r_data[41316] <= r_data[41315];
                
                r_data[41317] <= r_data[41316];
                
                r_data[41318] <= r_data[41317];
                
                r_data[41319] <= r_data[41318];
                
                r_data[41320] <= r_data[41319];
                
                r_data[41321] <= r_data[41320];
                
                r_data[41322] <= r_data[41321];
                
                r_data[41323] <= r_data[41322];
                
                r_data[41324] <= r_data[41323];
                
                r_data[41325] <= r_data[41324];
                
                r_data[41326] <= r_data[41325];
                
                r_data[41327] <= r_data[41326];
                
                r_data[41328] <= r_data[41327];
                
                r_data[41329] <= r_data[41328];
                
                r_data[41330] <= r_data[41329];
                
                r_data[41331] <= r_data[41330];
                
                r_data[41332] <= r_data[41331];
                
                r_data[41333] <= r_data[41332];
                
                r_data[41334] <= r_data[41333];
                
                r_data[41335] <= r_data[41334];
                
                r_data[41336] <= r_data[41335];
                
                r_data[41337] <= r_data[41336];
                
                r_data[41338] <= r_data[41337];
                
                r_data[41339] <= r_data[41338];
                
                r_data[41340] <= r_data[41339];
                
                r_data[41341] <= r_data[41340];
                
                r_data[41342] <= r_data[41341];
                
                r_data[41343] <= r_data[41342];
                
                r_data[41344] <= r_data[41343];
                
                r_data[41345] <= r_data[41344];
                
                r_data[41346] <= r_data[41345];
                
                r_data[41347] <= r_data[41346];
                
                r_data[41348] <= r_data[41347];
                
                r_data[41349] <= r_data[41348];
                
                r_data[41350] <= r_data[41349];
                
                r_data[41351] <= r_data[41350];
                
                r_data[41352] <= r_data[41351];
                
                r_data[41353] <= r_data[41352];
                
                r_data[41354] <= r_data[41353];
                
                r_data[41355] <= r_data[41354];
                
                r_data[41356] <= r_data[41355];
                
                r_data[41357] <= r_data[41356];
                
                r_data[41358] <= r_data[41357];
                
                r_data[41359] <= r_data[41358];
                
                r_data[41360] <= r_data[41359];
                
                r_data[41361] <= r_data[41360];
                
                r_data[41362] <= r_data[41361];
                
                r_data[41363] <= r_data[41362];
                
                r_data[41364] <= r_data[41363];
                
                r_data[41365] <= r_data[41364];
                
                r_data[41366] <= r_data[41365];
                
                r_data[41367] <= r_data[41366];
                
                r_data[41368] <= r_data[41367];
                
                r_data[41369] <= r_data[41368];
                
                r_data[41370] <= r_data[41369];
                
                r_data[41371] <= r_data[41370];
                
                r_data[41372] <= r_data[41371];
                
                r_data[41373] <= r_data[41372];
                
                r_data[41374] <= r_data[41373];
                
                r_data[41375] <= r_data[41374];
                
                r_data[41376] <= r_data[41375];
                
                r_data[41377] <= r_data[41376];
                
                r_data[41378] <= r_data[41377];
                
                r_data[41379] <= r_data[41378];
                
                r_data[41380] <= r_data[41379];
                
                r_data[41381] <= r_data[41380];
                
                r_data[41382] <= r_data[41381];
                
                r_data[41383] <= r_data[41382];
                
                r_data[41384] <= r_data[41383];
                
                r_data[41385] <= r_data[41384];
                
                r_data[41386] <= r_data[41385];
                
                r_data[41387] <= r_data[41386];
                
                r_data[41388] <= r_data[41387];
                
                r_data[41389] <= r_data[41388];
                
                r_data[41390] <= r_data[41389];
                
                r_data[41391] <= r_data[41390];
                
                r_data[41392] <= r_data[41391];
                
                r_data[41393] <= r_data[41392];
                
                r_data[41394] <= r_data[41393];
                
                r_data[41395] <= r_data[41394];
                
                r_data[41396] <= r_data[41395];
                
                r_data[41397] <= r_data[41396];
                
                r_data[41398] <= r_data[41397];
                
                r_data[41399] <= r_data[41398];
                
                r_data[41400] <= r_data[41399];
                
                r_data[41401] <= r_data[41400];
                
                r_data[41402] <= r_data[41401];
                
                r_data[41403] <= r_data[41402];
                
                r_data[41404] <= r_data[41403];
                
                r_data[41405] <= r_data[41404];
                
                r_data[41406] <= r_data[41405];
                
                r_data[41407] <= r_data[41406];
                
                r_data[41408] <= r_data[41407];
                
                r_data[41409] <= r_data[41408];
                
                r_data[41410] <= r_data[41409];
                
                r_data[41411] <= r_data[41410];
                
                r_data[41412] <= r_data[41411];
                
                r_data[41413] <= r_data[41412];
                
                r_data[41414] <= r_data[41413];
                
                r_data[41415] <= r_data[41414];
                
                r_data[41416] <= r_data[41415];
                
                r_data[41417] <= r_data[41416];
                
                r_data[41418] <= r_data[41417];
                
                r_data[41419] <= r_data[41418];
                
                r_data[41420] <= r_data[41419];
                
                r_data[41421] <= r_data[41420];
                
                r_data[41422] <= r_data[41421];
                
                r_data[41423] <= r_data[41422];
                
                r_data[41424] <= r_data[41423];
                
                r_data[41425] <= r_data[41424];
                
                r_data[41426] <= r_data[41425];
                
                r_data[41427] <= r_data[41426];
                
                r_data[41428] <= r_data[41427];
                
                r_data[41429] <= r_data[41428];
                
                r_data[41430] <= r_data[41429];
                
                r_data[41431] <= r_data[41430];
                
                r_data[41432] <= r_data[41431];
                
                r_data[41433] <= r_data[41432];
                
                r_data[41434] <= r_data[41433];
                
                r_data[41435] <= r_data[41434];
                
                r_data[41436] <= r_data[41435];
                
                r_data[41437] <= r_data[41436];
                
                r_data[41438] <= r_data[41437];
                
                r_data[41439] <= r_data[41438];
                
                r_data[41440] <= r_data[41439];
                
                r_data[41441] <= r_data[41440];
                
                r_data[41442] <= r_data[41441];
                
                r_data[41443] <= r_data[41442];
                
                r_data[41444] <= r_data[41443];
                
                r_data[41445] <= r_data[41444];
                
                r_data[41446] <= r_data[41445];
                
                r_data[41447] <= r_data[41446];
                
                r_data[41448] <= r_data[41447];
                
                r_data[41449] <= r_data[41448];
                
                r_data[41450] <= r_data[41449];
                
                r_data[41451] <= r_data[41450];
                
                r_data[41452] <= r_data[41451];
                
                r_data[41453] <= r_data[41452];
                
                r_data[41454] <= r_data[41453];
                
                r_data[41455] <= r_data[41454];
                
                r_data[41456] <= r_data[41455];
                
                r_data[41457] <= r_data[41456];
                
                r_data[41458] <= r_data[41457];
                
                r_data[41459] <= r_data[41458];
                
                r_data[41460] <= r_data[41459];
                
                r_data[41461] <= r_data[41460];
                
                r_data[41462] <= r_data[41461];
                
                r_data[41463] <= r_data[41462];
                
                r_data[41464] <= r_data[41463];
                
                r_data[41465] <= r_data[41464];
                
                r_data[41466] <= r_data[41465];
                
                r_data[41467] <= r_data[41466];
                
                r_data[41468] <= r_data[41467];
                
                r_data[41469] <= r_data[41468];
                
                r_data[41470] <= r_data[41469];
                
                r_data[41471] <= r_data[41470];
                
                r_data[41472] <= r_data[41471];
                
                r_data[41473] <= r_data[41472];
                
                r_data[41474] <= r_data[41473];
                
                r_data[41475] <= r_data[41474];
                
                r_data[41476] <= r_data[41475];
                
                r_data[41477] <= r_data[41476];
                
                r_data[41478] <= r_data[41477];
                
                r_data[41479] <= r_data[41478];
                
                r_data[41480] <= r_data[41479];
                
                r_data[41481] <= r_data[41480];
                
                r_data[41482] <= r_data[41481];
                
                r_data[41483] <= r_data[41482];
                
                r_data[41484] <= r_data[41483];
                
                r_data[41485] <= r_data[41484];
                
                r_data[41486] <= r_data[41485];
                
                r_data[41487] <= r_data[41486];
                
                r_data[41488] <= r_data[41487];
                
                r_data[41489] <= r_data[41488];
                
                r_data[41490] <= r_data[41489];
                
                r_data[41491] <= r_data[41490];
                
                r_data[41492] <= r_data[41491];
                
                r_data[41493] <= r_data[41492];
                
                r_data[41494] <= r_data[41493];
                
                r_data[41495] <= r_data[41494];
                
                r_data[41496] <= r_data[41495];
                
                r_data[41497] <= r_data[41496];
                
                r_data[41498] <= r_data[41497];
                
                r_data[41499] <= r_data[41498];
                
                r_data[41500] <= r_data[41499];
                
                r_data[41501] <= r_data[41500];
                
                r_data[41502] <= r_data[41501];
                
                r_data[41503] <= r_data[41502];
                
                r_data[41504] <= r_data[41503];
                
                r_data[41505] <= r_data[41504];
                
                r_data[41506] <= r_data[41505];
                
                r_data[41507] <= r_data[41506];
                
                r_data[41508] <= r_data[41507];
                
                r_data[41509] <= r_data[41508];
                
                r_data[41510] <= r_data[41509];
                
                r_data[41511] <= r_data[41510];
                
                r_data[41512] <= r_data[41511];
                
                r_data[41513] <= r_data[41512];
                
                r_data[41514] <= r_data[41513];
                
                r_data[41515] <= r_data[41514];
                
                r_data[41516] <= r_data[41515];
                
                r_data[41517] <= r_data[41516];
                
                r_data[41518] <= r_data[41517];
                
                r_data[41519] <= r_data[41518];
                
                r_data[41520] <= r_data[41519];
                
                r_data[41521] <= r_data[41520];
                
                r_data[41522] <= r_data[41521];
                
                r_data[41523] <= r_data[41522];
                
                r_data[41524] <= r_data[41523];
                
                r_data[41525] <= r_data[41524];
                
                r_data[41526] <= r_data[41525];
                
                r_data[41527] <= r_data[41526];
                
                r_data[41528] <= r_data[41527];
                
                r_data[41529] <= r_data[41528];
                
                r_data[41530] <= r_data[41529];
                
                r_data[41531] <= r_data[41530];
                
                r_data[41532] <= r_data[41531];
                
                r_data[41533] <= r_data[41532];
                
                r_data[41534] <= r_data[41533];
                
                r_data[41535] <= r_data[41534];
                
                r_data[41536] <= r_data[41535];
                
                r_data[41537] <= r_data[41536];
                
                r_data[41538] <= r_data[41537];
                
                r_data[41539] <= r_data[41538];
                
                r_data[41540] <= r_data[41539];
                
                r_data[41541] <= r_data[41540];
                
                r_data[41542] <= r_data[41541];
                
                r_data[41543] <= r_data[41542];
                
                r_data[41544] <= r_data[41543];
                
                r_data[41545] <= r_data[41544];
                
                r_data[41546] <= r_data[41545];
                
                r_data[41547] <= r_data[41546];
                
                r_data[41548] <= r_data[41547];
                
                r_data[41549] <= r_data[41548];
                
                r_data[41550] <= r_data[41549];
                
                r_data[41551] <= r_data[41550];
                
                r_data[41552] <= r_data[41551];
                
                r_data[41553] <= r_data[41552];
                
                r_data[41554] <= r_data[41553];
                
                r_data[41555] <= r_data[41554];
                
                r_data[41556] <= r_data[41555];
                
                r_data[41557] <= r_data[41556];
                
                r_data[41558] <= r_data[41557];
                
                r_data[41559] <= r_data[41558];
                
                r_data[41560] <= r_data[41559];
                
                r_data[41561] <= r_data[41560];
                
                r_data[41562] <= r_data[41561];
                
                r_data[41563] <= r_data[41562];
                
                r_data[41564] <= r_data[41563];
                
                r_data[41565] <= r_data[41564];
                
                r_data[41566] <= r_data[41565];
                
                r_data[41567] <= r_data[41566];
                
                r_data[41568] <= r_data[41567];
                
                r_data[41569] <= r_data[41568];
                
                r_data[41570] <= r_data[41569];
                
                r_data[41571] <= r_data[41570];
                
                r_data[41572] <= r_data[41571];
                
                r_data[41573] <= r_data[41572];
                
                r_data[41574] <= r_data[41573];
                
                r_data[41575] <= r_data[41574];
                
                r_data[41576] <= r_data[41575];
                
                r_data[41577] <= r_data[41576];
                
                r_data[41578] <= r_data[41577];
                
                r_data[41579] <= r_data[41578];
                
                r_data[41580] <= r_data[41579];
                
                r_data[41581] <= r_data[41580];
                
                r_data[41582] <= r_data[41581];
                
                r_data[41583] <= r_data[41582];
                
                r_data[41584] <= r_data[41583];
                
                r_data[41585] <= r_data[41584];
                
                r_data[41586] <= r_data[41585];
                
                r_data[41587] <= r_data[41586];
                
                r_data[41588] <= r_data[41587];
                
                r_data[41589] <= r_data[41588];
                
                r_data[41590] <= r_data[41589];
                
                r_data[41591] <= r_data[41590];
                
                r_data[41592] <= r_data[41591];
                
                r_data[41593] <= r_data[41592];
                
                r_data[41594] <= r_data[41593];
                
                r_data[41595] <= r_data[41594];
                
                r_data[41596] <= r_data[41595];
                
                r_data[41597] <= r_data[41596];
                
                r_data[41598] <= r_data[41597];
                
                r_data[41599] <= r_data[41598];
                
                r_data[41600] <= r_data[41599];
                
                r_data[41601] <= r_data[41600];
                
                r_data[41602] <= r_data[41601];
                
                r_data[41603] <= r_data[41602];
                
                r_data[41604] <= r_data[41603];
                
                r_data[41605] <= r_data[41604];
                
                r_data[41606] <= r_data[41605];
                
                r_data[41607] <= r_data[41606];
                
                r_data[41608] <= r_data[41607];
                
                r_data[41609] <= r_data[41608];
                
                r_data[41610] <= r_data[41609];
                
                r_data[41611] <= r_data[41610];
                
                r_data[41612] <= r_data[41611];
                
                r_data[41613] <= r_data[41612];
                
                r_data[41614] <= r_data[41613];
                
                r_data[41615] <= r_data[41614];
                
                r_data[41616] <= r_data[41615];
                
                r_data[41617] <= r_data[41616];
                
                r_data[41618] <= r_data[41617];
                
                r_data[41619] <= r_data[41618];
                
                r_data[41620] <= r_data[41619];
                
                r_data[41621] <= r_data[41620];
                
                r_data[41622] <= r_data[41621];
                
                r_data[41623] <= r_data[41622];
                
                r_data[41624] <= r_data[41623];
                
                r_data[41625] <= r_data[41624];
                
                r_data[41626] <= r_data[41625];
                
                r_data[41627] <= r_data[41626];
                
                r_data[41628] <= r_data[41627];
                
                r_data[41629] <= r_data[41628];
                
                r_data[41630] <= r_data[41629];
                
                r_data[41631] <= r_data[41630];
                
                r_data[41632] <= r_data[41631];
                
                r_data[41633] <= r_data[41632];
                
                r_data[41634] <= r_data[41633];
                
                r_data[41635] <= r_data[41634];
                
                r_data[41636] <= r_data[41635];
                
                r_data[41637] <= r_data[41636];
                
                r_data[41638] <= r_data[41637];
                
                r_data[41639] <= r_data[41638];
                
                r_data[41640] <= r_data[41639];
                
                r_data[41641] <= r_data[41640];
                
                r_data[41642] <= r_data[41641];
                
                r_data[41643] <= r_data[41642];
                
                r_data[41644] <= r_data[41643];
                
                r_data[41645] <= r_data[41644];
                
                r_data[41646] <= r_data[41645];
                
                r_data[41647] <= r_data[41646];
                
                r_data[41648] <= r_data[41647];
                
                r_data[41649] <= r_data[41648];
                
                r_data[41650] <= r_data[41649];
                
                r_data[41651] <= r_data[41650];
                
                r_data[41652] <= r_data[41651];
                
                r_data[41653] <= r_data[41652];
                
                r_data[41654] <= r_data[41653];
                
                r_data[41655] <= r_data[41654];
                
                r_data[41656] <= r_data[41655];
                
                r_data[41657] <= r_data[41656];
                
                r_data[41658] <= r_data[41657];
                
                r_data[41659] <= r_data[41658];
                
                r_data[41660] <= r_data[41659];
                
                r_data[41661] <= r_data[41660];
                
                r_data[41662] <= r_data[41661];
                
                r_data[41663] <= r_data[41662];
                
                r_data[41664] <= r_data[41663];
                
                r_data[41665] <= r_data[41664];
                
                r_data[41666] <= r_data[41665];
                
                r_data[41667] <= r_data[41666];
                
                r_data[41668] <= r_data[41667];
                
                r_data[41669] <= r_data[41668];
                
                r_data[41670] <= r_data[41669];
                
                r_data[41671] <= r_data[41670];
                
                r_data[41672] <= r_data[41671];
                
                r_data[41673] <= r_data[41672];
                
                r_data[41674] <= r_data[41673];
                
                r_data[41675] <= r_data[41674];
                
                r_data[41676] <= r_data[41675];
                
                r_data[41677] <= r_data[41676];
                
                r_data[41678] <= r_data[41677];
                
                r_data[41679] <= r_data[41678];
                
                r_data[41680] <= r_data[41679];
                
                r_data[41681] <= r_data[41680];
                
                r_data[41682] <= r_data[41681];
                
                r_data[41683] <= r_data[41682];
                
                r_data[41684] <= r_data[41683];
                
                r_data[41685] <= r_data[41684];
                
                r_data[41686] <= r_data[41685];
                
                r_data[41687] <= r_data[41686];
                
                r_data[41688] <= r_data[41687];
                
                r_data[41689] <= r_data[41688];
                
                r_data[41690] <= r_data[41689];
                
                r_data[41691] <= r_data[41690];
                
                r_data[41692] <= r_data[41691];
                
                r_data[41693] <= r_data[41692];
                
                r_data[41694] <= r_data[41693];
                
                r_data[41695] <= r_data[41694];
                
                r_data[41696] <= r_data[41695];
                
                r_data[41697] <= r_data[41696];
                
                r_data[41698] <= r_data[41697];
                
                r_data[41699] <= r_data[41698];
                
                r_data[41700] <= r_data[41699];
                
                r_data[41701] <= r_data[41700];
                
                r_data[41702] <= r_data[41701];
                
                r_data[41703] <= r_data[41702];
                
                r_data[41704] <= r_data[41703];
                
                r_data[41705] <= r_data[41704];
                
                r_data[41706] <= r_data[41705];
                
                r_data[41707] <= r_data[41706];
                
                r_data[41708] <= r_data[41707];
                
                r_data[41709] <= r_data[41708];
                
                r_data[41710] <= r_data[41709];
                
                r_data[41711] <= r_data[41710];
                
                r_data[41712] <= r_data[41711];
                
                r_data[41713] <= r_data[41712];
                
                r_data[41714] <= r_data[41713];
                
                r_data[41715] <= r_data[41714];
                
                r_data[41716] <= r_data[41715];
                
                r_data[41717] <= r_data[41716];
                
                r_data[41718] <= r_data[41717];
                
                r_data[41719] <= r_data[41718];
                
                r_data[41720] <= r_data[41719];
                
                r_data[41721] <= r_data[41720];
                
                r_data[41722] <= r_data[41721];
                
                r_data[41723] <= r_data[41722];
                
                r_data[41724] <= r_data[41723];
                
                r_data[41725] <= r_data[41724];
                
                r_data[41726] <= r_data[41725];
                
                r_data[41727] <= r_data[41726];
                
                r_data[41728] <= r_data[41727];
                
                r_data[41729] <= r_data[41728];
                
                r_data[41730] <= r_data[41729];
                
                r_data[41731] <= r_data[41730];
                
                r_data[41732] <= r_data[41731];
                
                r_data[41733] <= r_data[41732];
                
                r_data[41734] <= r_data[41733];
                
                r_data[41735] <= r_data[41734];
                
                r_data[41736] <= r_data[41735];
                
                r_data[41737] <= r_data[41736];
                
                r_data[41738] <= r_data[41737];
                
                r_data[41739] <= r_data[41738];
                
                r_data[41740] <= r_data[41739];
                
                r_data[41741] <= r_data[41740];
                
                r_data[41742] <= r_data[41741];
                
                r_data[41743] <= r_data[41742];
                
                r_data[41744] <= r_data[41743];
                
                r_data[41745] <= r_data[41744];
                
                r_data[41746] <= r_data[41745];
                
                r_data[41747] <= r_data[41746];
                
                r_data[41748] <= r_data[41747];
                
                r_data[41749] <= r_data[41748];
                
                r_data[41750] <= r_data[41749];
                
                r_data[41751] <= r_data[41750];
                
                r_data[41752] <= r_data[41751];
                
                r_data[41753] <= r_data[41752];
                
                r_data[41754] <= r_data[41753];
                
                r_data[41755] <= r_data[41754];
                
                r_data[41756] <= r_data[41755];
                
                r_data[41757] <= r_data[41756];
                
                r_data[41758] <= r_data[41757];
                
                r_data[41759] <= r_data[41758];
                
                r_data[41760] <= r_data[41759];
                
                r_data[41761] <= r_data[41760];
                
                r_data[41762] <= r_data[41761];
                
                r_data[41763] <= r_data[41762];
                
                r_data[41764] <= r_data[41763];
                
                r_data[41765] <= r_data[41764];
                
                r_data[41766] <= r_data[41765];
                
                r_data[41767] <= r_data[41766];
                
                r_data[41768] <= r_data[41767];
                
                r_data[41769] <= r_data[41768];
                
                r_data[41770] <= r_data[41769];
                
                r_data[41771] <= r_data[41770];
                
                r_data[41772] <= r_data[41771];
                
                r_data[41773] <= r_data[41772];
                
                r_data[41774] <= r_data[41773];
                
                r_data[41775] <= r_data[41774];
                
                r_data[41776] <= r_data[41775];
                
                r_data[41777] <= r_data[41776];
                
                r_data[41778] <= r_data[41777];
                
                r_data[41779] <= r_data[41778];
                
                r_data[41780] <= r_data[41779];
                
                r_data[41781] <= r_data[41780];
                
                r_data[41782] <= r_data[41781];
                
                r_data[41783] <= r_data[41782];
                
                r_data[41784] <= r_data[41783];
                
                r_data[41785] <= r_data[41784];
                
                r_data[41786] <= r_data[41785];
                
                r_data[41787] <= r_data[41786];
                
                r_data[41788] <= r_data[41787];
                
                r_data[41789] <= r_data[41788];
                
                r_data[41790] <= r_data[41789];
                
                r_data[41791] <= r_data[41790];
                
                r_data[41792] <= r_data[41791];
                
                r_data[41793] <= r_data[41792];
                
                r_data[41794] <= r_data[41793];
                
                r_data[41795] <= r_data[41794];
                
                r_data[41796] <= r_data[41795];
                
                r_data[41797] <= r_data[41796];
                
                r_data[41798] <= r_data[41797];
                
                r_data[41799] <= r_data[41798];
                
                r_data[41800] <= r_data[41799];
                
                r_data[41801] <= r_data[41800];
                
                r_data[41802] <= r_data[41801];
                
                r_data[41803] <= r_data[41802];
                
                r_data[41804] <= r_data[41803];
                
                r_data[41805] <= r_data[41804];
                
                r_data[41806] <= r_data[41805];
                
                r_data[41807] <= r_data[41806];
                
                r_data[41808] <= r_data[41807];
                
                r_data[41809] <= r_data[41808];
                
                r_data[41810] <= r_data[41809];
                
                r_data[41811] <= r_data[41810];
                
                r_data[41812] <= r_data[41811];
                
                r_data[41813] <= r_data[41812];
                
                r_data[41814] <= r_data[41813];
                
                r_data[41815] <= r_data[41814];
                
                r_data[41816] <= r_data[41815];
                
                r_data[41817] <= r_data[41816];
                
                r_data[41818] <= r_data[41817];
                
                r_data[41819] <= r_data[41818];
                
                r_data[41820] <= r_data[41819];
                
                r_data[41821] <= r_data[41820];
                
                r_data[41822] <= r_data[41821];
                
                r_data[41823] <= r_data[41822];
                
                r_data[41824] <= r_data[41823];
                
                r_data[41825] <= r_data[41824];
                
                r_data[41826] <= r_data[41825];
                
                r_data[41827] <= r_data[41826];
                
                r_data[41828] <= r_data[41827];
                
                r_data[41829] <= r_data[41828];
                
                r_data[41830] <= r_data[41829];
                
                r_data[41831] <= r_data[41830];
                
                r_data[41832] <= r_data[41831];
                
                r_data[41833] <= r_data[41832];
                
                r_data[41834] <= r_data[41833];
                
                r_data[41835] <= r_data[41834];
                
                r_data[41836] <= r_data[41835];
                
                r_data[41837] <= r_data[41836];
                
                r_data[41838] <= r_data[41837];
                
                r_data[41839] <= r_data[41838];
                
                r_data[41840] <= r_data[41839];
                
                r_data[41841] <= r_data[41840];
                
                r_data[41842] <= r_data[41841];
                
                r_data[41843] <= r_data[41842];
                
                r_data[41844] <= r_data[41843];
                
                r_data[41845] <= r_data[41844];
                
                r_data[41846] <= r_data[41845];
                
                r_data[41847] <= r_data[41846];
                
                r_data[41848] <= r_data[41847];
                
                r_data[41849] <= r_data[41848];
                
                r_data[41850] <= r_data[41849];
                
                r_data[41851] <= r_data[41850];
                
                r_data[41852] <= r_data[41851];
                
                r_data[41853] <= r_data[41852];
                
                r_data[41854] <= r_data[41853];
                
                r_data[41855] <= r_data[41854];
                
                r_data[41856] <= r_data[41855];
                
                r_data[41857] <= r_data[41856];
                
                r_data[41858] <= r_data[41857];
                
                r_data[41859] <= r_data[41858];
                
                r_data[41860] <= r_data[41859];
                
                r_data[41861] <= r_data[41860];
                
                r_data[41862] <= r_data[41861];
                
                r_data[41863] <= r_data[41862];
                
                r_data[41864] <= r_data[41863];
                
                r_data[41865] <= r_data[41864];
                
                r_data[41866] <= r_data[41865];
                
                r_data[41867] <= r_data[41866];
                
                r_data[41868] <= r_data[41867];
                
                r_data[41869] <= r_data[41868];
                
                r_data[41870] <= r_data[41869];
                
                r_data[41871] <= r_data[41870];
                
                r_data[41872] <= r_data[41871];
                
                r_data[41873] <= r_data[41872];
                
                r_data[41874] <= r_data[41873];
                
                r_data[41875] <= r_data[41874];
                
                r_data[41876] <= r_data[41875];
                
                r_data[41877] <= r_data[41876];
                
                r_data[41878] <= r_data[41877];
                
                r_data[41879] <= r_data[41878];
                
                r_data[41880] <= r_data[41879];
                
                r_data[41881] <= r_data[41880];
                
                r_data[41882] <= r_data[41881];
                
                r_data[41883] <= r_data[41882];
                
                r_data[41884] <= r_data[41883];
                
                r_data[41885] <= r_data[41884];
                
                r_data[41886] <= r_data[41885];
                
                r_data[41887] <= r_data[41886];
                
                r_data[41888] <= r_data[41887];
                
                r_data[41889] <= r_data[41888];
                
                r_data[41890] <= r_data[41889];
                
                r_data[41891] <= r_data[41890];
                
                r_data[41892] <= r_data[41891];
                
                r_data[41893] <= r_data[41892];
                
                r_data[41894] <= r_data[41893];
                
                r_data[41895] <= r_data[41894];
                
                r_data[41896] <= r_data[41895];
                
                r_data[41897] <= r_data[41896];
                
                r_data[41898] <= r_data[41897];
                
                r_data[41899] <= r_data[41898];
                
                r_data[41900] <= r_data[41899];
                
                r_data[41901] <= r_data[41900];
                
                r_data[41902] <= r_data[41901];
                
                r_data[41903] <= r_data[41902];
                
                r_data[41904] <= r_data[41903];
                
                r_data[41905] <= r_data[41904];
                
                r_data[41906] <= r_data[41905];
                
                r_data[41907] <= r_data[41906];
                
                r_data[41908] <= r_data[41907];
                
                r_data[41909] <= r_data[41908];
                
                r_data[41910] <= r_data[41909];
                
                r_data[41911] <= r_data[41910];
                
                r_data[41912] <= r_data[41911];
                
                r_data[41913] <= r_data[41912];
                
                r_data[41914] <= r_data[41913];
                
                r_data[41915] <= r_data[41914];
                
                r_data[41916] <= r_data[41915];
                
                r_data[41917] <= r_data[41916];
                
                r_data[41918] <= r_data[41917];
                
                r_data[41919] <= r_data[41918];
                
                r_data[41920] <= r_data[41919];
                
                r_data[41921] <= r_data[41920];
                
                r_data[41922] <= r_data[41921];
                
                r_data[41923] <= r_data[41922];
                
                r_data[41924] <= r_data[41923];
                
                r_data[41925] <= r_data[41924];
                
                r_data[41926] <= r_data[41925];
                
                r_data[41927] <= r_data[41926];
                
                r_data[41928] <= r_data[41927];
                
                r_data[41929] <= r_data[41928];
                
                r_data[41930] <= r_data[41929];
                
                r_data[41931] <= r_data[41930];
                
                r_data[41932] <= r_data[41931];
                
                r_data[41933] <= r_data[41932];
                
                r_data[41934] <= r_data[41933];
                
                r_data[41935] <= r_data[41934];
                
                r_data[41936] <= r_data[41935];
                
                r_data[41937] <= r_data[41936];
                
                r_data[41938] <= r_data[41937];
                
                r_data[41939] <= r_data[41938];
                
                r_data[41940] <= r_data[41939];
                
                r_data[41941] <= r_data[41940];
                
                r_data[41942] <= r_data[41941];
                
                r_data[41943] <= r_data[41942];
                
                r_data[41944] <= r_data[41943];
                
                r_data[41945] <= r_data[41944];
                
                r_data[41946] <= r_data[41945];
                
                r_data[41947] <= r_data[41946];
                
                r_data[41948] <= r_data[41947];
                
                r_data[41949] <= r_data[41948];
                
                r_data[41950] <= r_data[41949];
                
                r_data[41951] <= r_data[41950];
                
                r_data[41952] <= r_data[41951];
                
                r_data[41953] <= r_data[41952];
                
                r_data[41954] <= r_data[41953];
                
                r_data[41955] <= r_data[41954];
                
                r_data[41956] <= r_data[41955];
                
                r_data[41957] <= r_data[41956];
                
                r_data[41958] <= r_data[41957];
                
                r_data[41959] <= r_data[41958];
                
                r_data[41960] <= r_data[41959];
                
                r_data[41961] <= r_data[41960];
                
                r_data[41962] <= r_data[41961];
                
                r_data[41963] <= r_data[41962];
                
                r_data[41964] <= r_data[41963];
                
                r_data[41965] <= r_data[41964];
                
                r_data[41966] <= r_data[41965];
                
                r_data[41967] <= r_data[41966];
                
                r_data[41968] <= r_data[41967];
                
                r_data[41969] <= r_data[41968];
                
                r_data[41970] <= r_data[41969];
                
                r_data[41971] <= r_data[41970];
                
                r_data[41972] <= r_data[41971];
                
                r_data[41973] <= r_data[41972];
                
                r_data[41974] <= r_data[41973];
                
                r_data[41975] <= r_data[41974];
                
                r_data[41976] <= r_data[41975];
                
                r_data[41977] <= r_data[41976];
                
                r_data[41978] <= r_data[41977];
                
                r_data[41979] <= r_data[41978];
                
                r_data[41980] <= r_data[41979];
                
                r_data[41981] <= r_data[41980];
                
                r_data[41982] <= r_data[41981];
                
                r_data[41983] <= r_data[41982];
                
                r_data[41984] <= r_data[41983];
                
                r_data[41985] <= r_data[41984];
                
                r_data[41986] <= r_data[41985];
                
                r_data[41987] <= r_data[41986];
                
                r_data[41988] <= r_data[41987];
                
                r_data[41989] <= r_data[41988];
                
                r_data[41990] <= r_data[41989];
                
                r_data[41991] <= r_data[41990];
                
                r_data[41992] <= r_data[41991];
                
                r_data[41993] <= r_data[41992];
                
                r_data[41994] <= r_data[41993];
                
                r_data[41995] <= r_data[41994];
                
                r_data[41996] <= r_data[41995];
                
                r_data[41997] <= r_data[41996];
                
                r_data[41998] <= r_data[41997];
                
                r_data[41999] <= r_data[41998];
                
                r_data[42000] <= r_data[41999];
                
                r_data[42001] <= r_data[42000];
                
                r_data[42002] <= r_data[42001];
                
                r_data[42003] <= r_data[42002];
                
                r_data[42004] <= r_data[42003];
                
                r_data[42005] <= r_data[42004];
                
                r_data[42006] <= r_data[42005];
                
                r_data[42007] <= r_data[42006];
                
                r_data[42008] <= r_data[42007];
                
                r_data[42009] <= r_data[42008];
                
                r_data[42010] <= r_data[42009];
                
                r_data[42011] <= r_data[42010];
                
                r_data[42012] <= r_data[42011];
                
                r_data[42013] <= r_data[42012];
                
                r_data[42014] <= r_data[42013];
                
                r_data[42015] <= r_data[42014];
                
                r_data[42016] <= r_data[42015];
                
                r_data[42017] <= r_data[42016];
                
                r_data[42018] <= r_data[42017];
                
                r_data[42019] <= r_data[42018];
                
                r_data[42020] <= r_data[42019];
                
                r_data[42021] <= r_data[42020];
                
                r_data[42022] <= r_data[42021];
                
                r_data[42023] <= r_data[42022];
                
                r_data[42024] <= r_data[42023];
                
                r_data[42025] <= r_data[42024];
                
                r_data[42026] <= r_data[42025];
                
                r_data[42027] <= r_data[42026];
                
                r_data[42028] <= r_data[42027];
                
                r_data[42029] <= r_data[42028];
                
                r_data[42030] <= r_data[42029];
                
                r_data[42031] <= r_data[42030];
                
                r_data[42032] <= r_data[42031];
                
                r_data[42033] <= r_data[42032];
                
                r_data[42034] <= r_data[42033];
                
                r_data[42035] <= r_data[42034];
                
                r_data[42036] <= r_data[42035];
                
                r_data[42037] <= r_data[42036];
                
                r_data[42038] <= r_data[42037];
                
                r_data[42039] <= r_data[42038];
                
                r_data[42040] <= r_data[42039];
                
                r_data[42041] <= r_data[42040];
                
                r_data[42042] <= r_data[42041];
                
                r_data[42043] <= r_data[42042];
                
                r_data[42044] <= r_data[42043];
                
                r_data[42045] <= r_data[42044];
                
                r_data[42046] <= r_data[42045];
                
                r_data[42047] <= r_data[42046];
                
                r_data[42048] <= r_data[42047];
                
                r_data[42049] <= r_data[42048];
                
                r_data[42050] <= r_data[42049];
                
                r_data[42051] <= r_data[42050];
                
                r_data[42052] <= r_data[42051];
                
                r_data[42053] <= r_data[42052];
                
                r_data[42054] <= r_data[42053];
                
                r_data[42055] <= r_data[42054];
                
                r_data[42056] <= r_data[42055];
                
                r_data[42057] <= r_data[42056];
                
                r_data[42058] <= r_data[42057];
                
                r_data[42059] <= r_data[42058];
                
                r_data[42060] <= r_data[42059];
                
                r_data[42061] <= r_data[42060];
                
                r_data[42062] <= r_data[42061];
                
                r_data[42063] <= r_data[42062];
                
                r_data[42064] <= r_data[42063];
                
                r_data[42065] <= r_data[42064];
                
                r_data[42066] <= r_data[42065];
                
                r_data[42067] <= r_data[42066];
                
                r_data[42068] <= r_data[42067];
                
                r_data[42069] <= r_data[42068];
                
                r_data[42070] <= r_data[42069];
                
                r_data[42071] <= r_data[42070];
                
                r_data[42072] <= r_data[42071];
                
                r_data[42073] <= r_data[42072];
                
                r_data[42074] <= r_data[42073];
                
                r_data[42075] <= r_data[42074];
                
                r_data[42076] <= r_data[42075];
                
                r_data[42077] <= r_data[42076];
                
                r_data[42078] <= r_data[42077];
                
                r_data[42079] <= r_data[42078];
                
                r_data[42080] <= r_data[42079];
                
                r_data[42081] <= r_data[42080];
                
                r_data[42082] <= r_data[42081];
                
                r_data[42083] <= r_data[42082];
                
                r_data[42084] <= r_data[42083];
                
                r_data[42085] <= r_data[42084];
                
                r_data[42086] <= r_data[42085];
                
                r_data[42087] <= r_data[42086];
                
                r_data[42088] <= r_data[42087];
                
                r_data[42089] <= r_data[42088];
                
                r_data[42090] <= r_data[42089];
                
                r_data[42091] <= r_data[42090];
                
                r_data[42092] <= r_data[42091];
                
                r_data[42093] <= r_data[42092];
                
                r_data[42094] <= r_data[42093];
                
                r_data[42095] <= r_data[42094];
                
                r_data[42096] <= r_data[42095];
                
                r_data[42097] <= r_data[42096];
                
                r_data[42098] <= r_data[42097];
                
                r_data[42099] <= r_data[42098];
                
                r_data[42100] <= r_data[42099];
                
                r_data[42101] <= r_data[42100];
                
                r_data[42102] <= r_data[42101];
                
                r_data[42103] <= r_data[42102];
                
                r_data[42104] <= r_data[42103];
                
                r_data[42105] <= r_data[42104];
                
                r_data[42106] <= r_data[42105];
                
                r_data[42107] <= r_data[42106];
                
                r_data[42108] <= r_data[42107];
                
                r_data[42109] <= r_data[42108];
                
                r_data[42110] <= r_data[42109];
                
                r_data[42111] <= r_data[42110];
                
                r_data[42112] <= r_data[42111];
                
                r_data[42113] <= r_data[42112];
                
                r_data[42114] <= r_data[42113];
                
                r_data[42115] <= r_data[42114];
                
                r_data[42116] <= r_data[42115];
                
                r_data[42117] <= r_data[42116];
                
                r_data[42118] <= r_data[42117];
                
                r_data[42119] <= r_data[42118];
                
                r_data[42120] <= r_data[42119];
                
                r_data[42121] <= r_data[42120];
                
                r_data[42122] <= r_data[42121];
                
                r_data[42123] <= r_data[42122];
                
                r_data[42124] <= r_data[42123];
                
                r_data[42125] <= r_data[42124];
                
                r_data[42126] <= r_data[42125];
                
                r_data[42127] <= r_data[42126];
                
                r_data[42128] <= r_data[42127];
                
                r_data[42129] <= r_data[42128];
                
                r_data[42130] <= r_data[42129];
                
                r_data[42131] <= r_data[42130];
                
                r_data[42132] <= r_data[42131];
                
                r_data[42133] <= r_data[42132];
                
                r_data[42134] <= r_data[42133];
                
                r_data[42135] <= r_data[42134];
                
                r_data[42136] <= r_data[42135];
                
                r_data[42137] <= r_data[42136];
                
                r_data[42138] <= r_data[42137];
                
                r_data[42139] <= r_data[42138];
                
                r_data[42140] <= r_data[42139];
                
                r_data[42141] <= r_data[42140];
                
                r_data[42142] <= r_data[42141];
                
                r_data[42143] <= r_data[42142];
                
                r_data[42144] <= r_data[42143];
                
                r_data[42145] <= r_data[42144];
                
                r_data[42146] <= r_data[42145];
                
                r_data[42147] <= r_data[42146];
                
                r_data[42148] <= r_data[42147];
                
                r_data[42149] <= r_data[42148];
                
                r_data[42150] <= r_data[42149];
                
                r_data[42151] <= r_data[42150];
                
                r_data[42152] <= r_data[42151];
                
                r_data[42153] <= r_data[42152];
                
                r_data[42154] <= r_data[42153];
                
                r_data[42155] <= r_data[42154];
                
                r_data[42156] <= r_data[42155];
                
                r_data[42157] <= r_data[42156];
                
                r_data[42158] <= r_data[42157];
                
                r_data[42159] <= r_data[42158];
                
                r_data[42160] <= r_data[42159];
                
                r_data[42161] <= r_data[42160];
                
                r_data[42162] <= r_data[42161];
                
                r_data[42163] <= r_data[42162];
                
                r_data[42164] <= r_data[42163];
                
                r_data[42165] <= r_data[42164];
                
                r_data[42166] <= r_data[42165];
                
                r_data[42167] <= r_data[42166];
                
                r_data[42168] <= r_data[42167];
                
                r_data[42169] <= r_data[42168];
                
                r_data[42170] <= r_data[42169];
                
                r_data[42171] <= r_data[42170];
                
                r_data[42172] <= r_data[42171];
                
                r_data[42173] <= r_data[42172];
                
                r_data[42174] <= r_data[42173];
                
                r_data[42175] <= r_data[42174];
                
                r_data[42176] <= r_data[42175];
                
                r_data[42177] <= r_data[42176];
                
                r_data[42178] <= r_data[42177];
                
                r_data[42179] <= r_data[42178];
                
                r_data[42180] <= r_data[42179];
                
                r_data[42181] <= r_data[42180];
                
                r_data[42182] <= r_data[42181];
                
                r_data[42183] <= r_data[42182];
                
                r_data[42184] <= r_data[42183];
                
                r_data[42185] <= r_data[42184];
                
                r_data[42186] <= r_data[42185];
                
                r_data[42187] <= r_data[42186];
                
                r_data[42188] <= r_data[42187];
                
                r_data[42189] <= r_data[42188];
                
                r_data[42190] <= r_data[42189];
                
                r_data[42191] <= r_data[42190];
                
                r_data[42192] <= r_data[42191];
                
                r_data[42193] <= r_data[42192];
                
                r_data[42194] <= r_data[42193];
                
                r_data[42195] <= r_data[42194];
                
                r_data[42196] <= r_data[42195];
                
                r_data[42197] <= r_data[42196];
                
                r_data[42198] <= r_data[42197];
                
                r_data[42199] <= r_data[42198];
                
                r_data[42200] <= r_data[42199];
                
                r_data[42201] <= r_data[42200];
                
                r_data[42202] <= r_data[42201];
                
                r_data[42203] <= r_data[42202];
                
                r_data[42204] <= r_data[42203];
                
                r_data[42205] <= r_data[42204];
                
                r_data[42206] <= r_data[42205];
                
                r_data[42207] <= r_data[42206];
                
                r_data[42208] <= r_data[42207];
                
                r_data[42209] <= r_data[42208];
                
                r_data[42210] <= r_data[42209];
                
                r_data[42211] <= r_data[42210];
                
                r_data[42212] <= r_data[42211];
                
                r_data[42213] <= r_data[42212];
                
                r_data[42214] <= r_data[42213];
                
                r_data[42215] <= r_data[42214];
                
                r_data[42216] <= r_data[42215];
                
                r_data[42217] <= r_data[42216];
                
                r_data[42218] <= r_data[42217];
                
                r_data[42219] <= r_data[42218];
                
                r_data[42220] <= r_data[42219];
                
                r_data[42221] <= r_data[42220];
                
                r_data[42222] <= r_data[42221];
                
                r_data[42223] <= r_data[42222];
                
                r_data[42224] <= r_data[42223];
                
                r_data[42225] <= r_data[42224];
                
                r_data[42226] <= r_data[42225];
                
                r_data[42227] <= r_data[42226];
                
                r_data[42228] <= r_data[42227];
                
                r_data[42229] <= r_data[42228];
                
                r_data[42230] <= r_data[42229];
                
                r_data[42231] <= r_data[42230];
                
                r_data[42232] <= r_data[42231];
                
                r_data[42233] <= r_data[42232];
                
                r_data[42234] <= r_data[42233];
                
                r_data[42235] <= r_data[42234];
                
                r_data[42236] <= r_data[42235];
                
                r_data[42237] <= r_data[42236];
                
                r_data[42238] <= r_data[42237];
                
                r_data[42239] <= r_data[42238];
                
                r_data[42240] <= r_data[42239];
                
                r_data[42241] <= r_data[42240];
                
                r_data[42242] <= r_data[42241];
                
                r_data[42243] <= r_data[42242];
                
                r_data[42244] <= r_data[42243];
                
                r_data[42245] <= r_data[42244];
                
                r_data[42246] <= r_data[42245];
                
                r_data[42247] <= r_data[42246];
                
                r_data[42248] <= r_data[42247];
                
                r_data[42249] <= r_data[42248];
                
                r_data[42250] <= r_data[42249];
                
                r_data[42251] <= r_data[42250];
                
                r_data[42252] <= r_data[42251];
                
                r_data[42253] <= r_data[42252];
                
                r_data[42254] <= r_data[42253];
                
                r_data[42255] <= r_data[42254];
                
                r_data[42256] <= r_data[42255];
                
                r_data[42257] <= r_data[42256];
                
                r_data[42258] <= r_data[42257];
                
                r_data[42259] <= r_data[42258];
                
                r_data[42260] <= r_data[42259];
                
                r_data[42261] <= r_data[42260];
                
                r_data[42262] <= r_data[42261];
                
                r_data[42263] <= r_data[42262];
                
                r_data[42264] <= r_data[42263];
                
                r_data[42265] <= r_data[42264];
                
                r_data[42266] <= r_data[42265];
                
                r_data[42267] <= r_data[42266];
                
                r_data[42268] <= r_data[42267];
                
                r_data[42269] <= r_data[42268];
                
                r_data[42270] <= r_data[42269];
                
                r_data[42271] <= r_data[42270];
                
                r_data[42272] <= r_data[42271];
                
                r_data[42273] <= r_data[42272];
                
                r_data[42274] <= r_data[42273];
                
                r_data[42275] <= r_data[42274];
                
                r_data[42276] <= r_data[42275];
                
                r_data[42277] <= r_data[42276];
                
                r_data[42278] <= r_data[42277];
                
                r_data[42279] <= r_data[42278];
                
                r_data[42280] <= r_data[42279];
                
                r_data[42281] <= r_data[42280];
                
                r_data[42282] <= r_data[42281];
                
                r_data[42283] <= r_data[42282];
                
                r_data[42284] <= r_data[42283];
                
                r_data[42285] <= r_data[42284];
                
                r_data[42286] <= r_data[42285];
                
                r_data[42287] <= r_data[42286];
                
                r_data[42288] <= r_data[42287];
                
                r_data[42289] <= r_data[42288];
                
                r_data[42290] <= r_data[42289];
                
                r_data[42291] <= r_data[42290];
                
                r_data[42292] <= r_data[42291];
                
                r_data[42293] <= r_data[42292];
                
                r_data[42294] <= r_data[42293];
                
                r_data[42295] <= r_data[42294];
                
                r_data[42296] <= r_data[42295];
                
                r_data[42297] <= r_data[42296];
                
                r_data[42298] <= r_data[42297];
                
                r_data[42299] <= r_data[42298];
                
                r_data[42300] <= r_data[42299];
                
                r_data[42301] <= r_data[42300];
                
                r_data[42302] <= r_data[42301];
                
                r_data[42303] <= r_data[42302];
                
                r_data[42304] <= r_data[42303];
                
                r_data[42305] <= r_data[42304];
                
                r_data[42306] <= r_data[42305];
                
                r_data[42307] <= r_data[42306];
                
                r_data[42308] <= r_data[42307];
                
                r_data[42309] <= r_data[42308];
                
                r_data[42310] <= r_data[42309];
                
                r_data[42311] <= r_data[42310];
                
                r_data[42312] <= r_data[42311];
                
                r_data[42313] <= r_data[42312];
                
                r_data[42314] <= r_data[42313];
                
                r_data[42315] <= r_data[42314];
                
                r_data[42316] <= r_data[42315];
                
                r_data[42317] <= r_data[42316];
                
                r_data[42318] <= r_data[42317];
                
                r_data[42319] <= r_data[42318];
                
                r_data[42320] <= r_data[42319];
                
                r_data[42321] <= r_data[42320];
                
                r_data[42322] <= r_data[42321];
                
                r_data[42323] <= r_data[42322];
                
                r_data[42324] <= r_data[42323];
                
                r_data[42325] <= r_data[42324];
                
                r_data[42326] <= r_data[42325];
                
                r_data[42327] <= r_data[42326];
                
                r_data[42328] <= r_data[42327];
                
                r_data[42329] <= r_data[42328];
                
                r_data[42330] <= r_data[42329];
                
                r_data[42331] <= r_data[42330];
                
                r_data[42332] <= r_data[42331];
                
                r_data[42333] <= r_data[42332];
                
                r_data[42334] <= r_data[42333];
                
                r_data[42335] <= r_data[42334];
                
                r_data[42336] <= r_data[42335];
                
                r_data[42337] <= r_data[42336];
                
                r_data[42338] <= r_data[42337];
                
                r_data[42339] <= r_data[42338];
                
                r_data[42340] <= r_data[42339];
                
                r_data[42341] <= r_data[42340];
                
                r_data[42342] <= r_data[42341];
                
                r_data[42343] <= r_data[42342];
                
                r_data[42344] <= r_data[42343];
                
                r_data[42345] <= r_data[42344];
                
                r_data[42346] <= r_data[42345];
                
                r_data[42347] <= r_data[42346];
                
                r_data[42348] <= r_data[42347];
                
                r_data[42349] <= r_data[42348];
                
                r_data[42350] <= r_data[42349];
                
                r_data[42351] <= r_data[42350];
                
                r_data[42352] <= r_data[42351];
                
                r_data[42353] <= r_data[42352];
                
                r_data[42354] <= r_data[42353];
                
                r_data[42355] <= r_data[42354];
                
                r_data[42356] <= r_data[42355];
                
                r_data[42357] <= r_data[42356];
                
                r_data[42358] <= r_data[42357];
                
                r_data[42359] <= r_data[42358];
                
                r_data[42360] <= r_data[42359];
                
                r_data[42361] <= r_data[42360];
                
                r_data[42362] <= r_data[42361];
                
                r_data[42363] <= r_data[42362];
                
                r_data[42364] <= r_data[42363];
                
                r_data[42365] <= r_data[42364];
                
                r_data[42366] <= r_data[42365];
                
                r_data[42367] <= r_data[42366];
                
            end
        end
    end
    assign data_out = r_data;   

endmodule